-------------------------------------------------------------------------------
--
-- Final examination - Digital Logic Design
-- Alberto Boffi - Politecnico di Milano, AY 2020/21
-- TEST MODULE: Shift level = 5
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity shlev5_tb is
end shlev5_tb;

architecture shlev5tb of shlev5_tb is
constant c_CLOCK_PERIOD         : time := 15 ns;
signal   tb_done                : std_logic;
signal   mem_address            : std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst                 : std_logic := '0';
signal   tb_start               : std_logic := '0';
signal   tb_clk                 : std_logic := '0';
signal   mem_o_data,mem_i_data  : std_logic_vector (7 downto 0);
signal   enable_wire            : std_logic;
signal   mem_we                 : std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);


signal RAM: ram_type :=
	(0 => std_logic_vector(to_unsigned(59, 8)),
	1 => std_logic_vector(to_unsigned(71, 8)),
	2 => std_logic_vector(to_unsigned(171, 8)),
	3 => std_logic_vector(to_unsigned(173, 8)),
	4 => std_logic_vector(to_unsigned(170, 8)),
	5 => std_logic_vector(to_unsigned(164, 8)),
	6 => std_logic_vector(to_unsigned(168, 8)),
	7 => std_logic_vector(to_unsigned(170, 8)),
	8 => std_logic_vector(to_unsigned(169, 8)),
	9 => std_logic_vector(to_unsigned(165, 8)),
	10 => std_logic_vector(to_unsigned(163, 8)),
	11 => std_logic_vector(to_unsigned(169, 8)),
	12 => std_logic_vector(to_unsigned(164, 8)),
	13 => std_logic_vector(to_unsigned(170, 8)),
	14 => std_logic_vector(to_unsigned(172, 8)),
	15 => std_logic_vector(to_unsigned(166, 8)),
	16 => std_logic_vector(to_unsigned(162, 8)),
	17 => std_logic_vector(to_unsigned(164, 8)),
	18 => std_logic_vector(to_unsigned(171, 8)),
	19 => std_logic_vector(to_unsigned(171, 8)),
	20 => std_logic_vector(to_unsigned(173, 8)),
	21 => std_logic_vector(to_unsigned(176, 8)),
	22 => std_logic_vector(to_unsigned(169, 8)),
	23 => std_logic_vector(to_unsigned(174, 8)),
	24 => std_logic_vector(to_unsigned(167, 8)),
	25 => std_logic_vector(to_unsigned(174, 8)),
	26 => std_logic_vector(to_unsigned(170, 8)),
	27 => std_logic_vector(to_unsigned(169, 8)),
	28 => std_logic_vector(to_unsigned(170, 8)),
	29 => std_logic_vector(to_unsigned(165, 8)),
	30 => std_logic_vector(to_unsigned(172, 8)),
	31 => std_logic_vector(to_unsigned(163, 8)),
	32 => std_logic_vector(to_unsigned(173, 8)),
	33 => std_logic_vector(to_unsigned(170, 8)),
	34 => std_logic_vector(to_unsigned(169, 8)),
	35 => std_logic_vector(to_unsigned(169, 8)),
	36 => std_logic_vector(to_unsigned(162, 8)),
	37 => std_logic_vector(to_unsigned(175, 8)),
	38 => std_logic_vector(to_unsigned(176, 8)),
	39 => std_logic_vector(to_unsigned(176, 8)),
	40 => std_logic_vector(to_unsigned(169, 8)),
	41 => std_logic_vector(to_unsigned(174, 8)),
	42 => std_logic_vector(to_unsigned(162, 8)),
	43 => std_logic_vector(to_unsigned(168, 8)),
	44 => std_logic_vector(to_unsigned(162, 8)),
	45 => std_logic_vector(to_unsigned(164, 8)),
	46 => std_logic_vector(to_unsigned(162, 8)),
	47 => std_logic_vector(to_unsigned(169, 8)),
	48 => std_logic_vector(to_unsigned(166, 8)),
	49 => std_logic_vector(to_unsigned(162, 8)),
	50 => std_logic_vector(to_unsigned(166, 8)),
	51 => std_logic_vector(to_unsigned(170, 8)),
	52 => std_logic_vector(to_unsigned(164, 8)),
	53 => std_logic_vector(to_unsigned(168, 8)),
	54 => std_logic_vector(to_unsigned(164, 8)),
	55 => std_logic_vector(to_unsigned(173, 8)),
	56 => std_logic_vector(to_unsigned(167, 8)),
	57 => std_logic_vector(to_unsigned(166, 8)),
	58 => std_logic_vector(to_unsigned(169, 8)),
	59 => std_logic_vector(to_unsigned(167, 8)),
	60 => std_logic_vector(to_unsigned(168, 8)),
	61 => std_logic_vector(to_unsigned(171, 8)),
	62 => std_logic_vector(to_unsigned(167, 8)),
	63 => std_logic_vector(to_unsigned(162, 8)),
	64 => std_logic_vector(to_unsigned(167, 8)),
	65 => std_logic_vector(to_unsigned(166, 8)),
	66 => std_logic_vector(to_unsigned(171, 8)),
	67 => std_logic_vector(to_unsigned(162, 8)),
	68 => std_logic_vector(to_unsigned(173, 8)),
	69 => std_logic_vector(to_unsigned(162, 8)),
	70 => std_logic_vector(to_unsigned(166, 8)),
	71 => std_logic_vector(to_unsigned(173, 8)),
	72 => std_logic_vector(to_unsigned(170, 8)),
	73 => std_logic_vector(to_unsigned(174, 8)),
	74 => std_logic_vector(to_unsigned(172, 8)),
	75 => std_logic_vector(to_unsigned(175, 8)),
	76 => std_logic_vector(to_unsigned(164, 8)),
	77 => std_logic_vector(to_unsigned(171, 8)),
	78 => std_logic_vector(to_unsigned(176, 8)),
	79 => std_logic_vector(to_unsigned(175, 8)),
	80 => std_logic_vector(to_unsigned(169, 8)),
	81 => std_logic_vector(to_unsigned(170, 8)),
	82 => std_logic_vector(to_unsigned(165, 8)),
	83 => std_logic_vector(to_unsigned(176, 8)),
	84 => std_logic_vector(to_unsigned(168, 8)),
	85 => std_logic_vector(to_unsigned(168, 8)),
	86 => std_logic_vector(to_unsigned(173, 8)),
	87 => std_logic_vector(to_unsigned(171, 8)),
	88 => std_logic_vector(to_unsigned(163, 8)),
	89 => std_logic_vector(to_unsigned(175, 8)),
	90 => std_logic_vector(to_unsigned(168, 8)),
	91 => std_logic_vector(to_unsigned(170, 8)),
	92 => std_logic_vector(to_unsigned(163, 8)),
	93 => std_logic_vector(to_unsigned(167, 8)),
	94 => std_logic_vector(to_unsigned(175, 8)),
	95 => std_logic_vector(to_unsigned(165, 8)),
	96 => std_logic_vector(to_unsigned(165, 8)),
	97 => std_logic_vector(to_unsigned(162, 8)),
	98 => std_logic_vector(to_unsigned(166, 8)),
	99 => std_logic_vector(to_unsigned(176, 8)),
	100 => std_logic_vector(to_unsigned(175, 8)),
	101 => std_logic_vector(to_unsigned(167, 8)),
	102 => std_logic_vector(to_unsigned(175, 8)),
	103 => std_logic_vector(to_unsigned(162, 8)),
	104 => std_logic_vector(to_unsigned(162, 8)),
	105 => std_logic_vector(to_unsigned(165, 8)),
	106 => std_logic_vector(to_unsigned(176, 8)),
	107 => std_logic_vector(to_unsigned(168, 8)),
	108 => std_logic_vector(to_unsigned(175, 8)),
	109 => std_logic_vector(to_unsigned(168, 8)),
	110 => std_logic_vector(to_unsigned(169, 8)),
	111 => std_logic_vector(to_unsigned(174, 8)),
	112 => std_logic_vector(to_unsigned(173, 8)),
	113 => std_logic_vector(to_unsigned(166, 8)),
	114 => std_logic_vector(to_unsigned(176, 8)),
	115 => std_logic_vector(to_unsigned(176, 8)),
	116 => std_logic_vector(to_unsigned(162, 8)),
	117 => std_logic_vector(to_unsigned(167, 8)),
	118 => std_logic_vector(to_unsigned(165, 8)),
	119 => std_logic_vector(to_unsigned(166, 8)),
	120 => std_logic_vector(to_unsigned(165, 8)),
	121 => std_logic_vector(to_unsigned(171, 8)),
	122 => std_logic_vector(to_unsigned(168, 8)),
	123 => std_logic_vector(to_unsigned(164, 8)),
	124 => std_logic_vector(to_unsigned(163, 8)),
	125 => std_logic_vector(to_unsigned(169, 8)),
	126 => std_logic_vector(to_unsigned(166, 8)),
	127 => std_logic_vector(to_unsigned(171, 8)),
	128 => std_logic_vector(to_unsigned(167, 8)),
	129 => std_logic_vector(to_unsigned(165, 8)),
	130 => std_logic_vector(to_unsigned(174, 8)),
	131 => std_logic_vector(to_unsigned(167, 8)),
	132 => std_logic_vector(to_unsigned(167, 8)),
	133 => std_logic_vector(to_unsigned(162, 8)),
	134 => std_logic_vector(to_unsigned(163, 8)),
	135 => std_logic_vector(to_unsigned(175, 8)),
	136 => std_logic_vector(to_unsigned(165, 8)),
	137 => std_logic_vector(to_unsigned(176, 8)),
	138 => std_logic_vector(to_unsigned(170, 8)),
	139 => std_logic_vector(to_unsigned(163, 8)),
	140 => std_logic_vector(to_unsigned(169, 8)),
	141 => std_logic_vector(to_unsigned(163, 8)),
	142 => std_logic_vector(to_unsigned(171, 8)),
	143 => std_logic_vector(to_unsigned(164, 8)),
	144 => std_logic_vector(to_unsigned(167, 8)),
	145 => std_logic_vector(to_unsigned(171, 8)),
	146 => std_logic_vector(to_unsigned(166, 8)),
	147 => std_logic_vector(to_unsigned(175, 8)),
	148 => std_logic_vector(to_unsigned(176, 8)),
	149 => std_logic_vector(to_unsigned(175, 8)),
	150 => std_logic_vector(to_unsigned(167, 8)),
	151 => std_logic_vector(to_unsigned(162, 8)),
	152 => std_logic_vector(to_unsigned(163, 8)),
	153 => std_logic_vector(to_unsigned(166, 8)),
	154 => std_logic_vector(to_unsigned(170, 8)),
	155 => std_logic_vector(to_unsigned(163, 8)),
	156 => std_logic_vector(to_unsigned(174, 8)),
	157 => std_logic_vector(to_unsigned(167, 8)),
	158 => std_logic_vector(to_unsigned(166, 8)),
	159 => std_logic_vector(to_unsigned(166, 8)),
	160 => std_logic_vector(to_unsigned(163, 8)),
	161 => std_logic_vector(to_unsigned(174, 8)),
	162 => std_logic_vector(to_unsigned(176, 8)),
	163 => std_logic_vector(to_unsigned(166, 8)),
	164 => std_logic_vector(to_unsigned(172, 8)),
	165 => std_logic_vector(to_unsigned(165, 8)),
	166 => std_logic_vector(to_unsigned(170, 8)),
	167 => std_logic_vector(to_unsigned(170, 8)),
	168 => std_logic_vector(to_unsigned(168, 8)),
	169 => std_logic_vector(to_unsigned(171, 8)),
	170 => std_logic_vector(to_unsigned(164, 8)),
	171 => std_logic_vector(to_unsigned(163, 8)),
	172 => std_logic_vector(to_unsigned(171, 8)),
	173 => std_logic_vector(to_unsigned(173, 8)),
	174 => std_logic_vector(to_unsigned(168, 8)),
	175 => std_logic_vector(to_unsigned(167, 8)),
	176 => std_logic_vector(to_unsigned(162, 8)),
	177 => std_logic_vector(to_unsigned(174, 8)),
	178 => std_logic_vector(to_unsigned(163, 8)),
	179 => std_logic_vector(to_unsigned(171, 8)),
	180 => std_logic_vector(to_unsigned(166, 8)),
	181 => std_logic_vector(to_unsigned(169, 8)),
	182 => std_logic_vector(to_unsigned(171, 8)),
	183 => std_logic_vector(to_unsigned(170, 8)),
	184 => std_logic_vector(to_unsigned(169, 8)),
	185 => std_logic_vector(to_unsigned(162, 8)),
	186 => std_logic_vector(to_unsigned(170, 8)),
	187 => std_logic_vector(to_unsigned(171, 8)),
	188 => std_logic_vector(to_unsigned(169, 8)),
	189 => std_logic_vector(to_unsigned(167, 8)),
	190 => std_logic_vector(to_unsigned(164, 8)),
	191 => std_logic_vector(to_unsigned(175, 8)),
	192 => std_logic_vector(to_unsigned(172, 8)),
	193 => std_logic_vector(to_unsigned(169, 8)),
	194 => std_logic_vector(to_unsigned(163, 8)),
	195 => std_logic_vector(to_unsigned(162, 8)),
	196 => std_logic_vector(to_unsigned(162, 8)),
	197 => std_logic_vector(to_unsigned(169, 8)),
	198 => std_logic_vector(to_unsigned(173, 8)),
	199 => std_logic_vector(to_unsigned(170, 8)),
	200 => std_logic_vector(to_unsigned(162, 8)),
	201 => std_logic_vector(to_unsigned(166, 8)),
	202 => std_logic_vector(to_unsigned(165, 8)),
	203 => std_logic_vector(to_unsigned(168, 8)),
	204 => std_logic_vector(to_unsigned(165, 8)),
	205 => std_logic_vector(to_unsigned(175, 8)),
	206 => std_logic_vector(to_unsigned(164, 8)),
	207 => std_logic_vector(to_unsigned(164, 8)),
	208 => std_logic_vector(to_unsigned(174, 8)),
	209 => std_logic_vector(to_unsigned(172, 8)),
	210 => std_logic_vector(to_unsigned(174, 8)),
	211 => std_logic_vector(to_unsigned(171, 8)),
	212 => std_logic_vector(to_unsigned(173, 8)),
	213 => std_logic_vector(to_unsigned(167, 8)),
	214 => std_logic_vector(to_unsigned(166, 8)),
	215 => std_logic_vector(to_unsigned(168, 8)),
	216 => std_logic_vector(to_unsigned(168, 8)),
	217 => std_logic_vector(to_unsigned(168, 8)),
	218 => std_logic_vector(to_unsigned(163, 8)),
	219 => std_logic_vector(to_unsigned(173, 8)),
	220 => std_logic_vector(to_unsigned(169, 8)),
	221 => std_logic_vector(to_unsigned(169, 8)),
	222 => std_logic_vector(to_unsigned(164, 8)),
	223 => std_logic_vector(to_unsigned(168, 8)),
	224 => std_logic_vector(to_unsigned(171, 8)),
	225 => std_logic_vector(to_unsigned(163, 8)),
	226 => std_logic_vector(to_unsigned(168, 8)),
	227 => std_logic_vector(to_unsigned(174, 8)),
	228 => std_logic_vector(to_unsigned(170, 8)),
	229 => std_logic_vector(to_unsigned(170, 8)),
	230 => std_logic_vector(to_unsigned(168, 8)),
	231 => std_logic_vector(to_unsigned(176, 8)),
	232 => std_logic_vector(to_unsigned(163, 8)),
	233 => std_logic_vector(to_unsigned(173, 8)),
	234 => std_logic_vector(to_unsigned(173, 8)),
	235 => std_logic_vector(to_unsigned(165, 8)),
	236 => std_logic_vector(to_unsigned(168, 8)),
	237 => std_logic_vector(to_unsigned(168, 8)),
	238 => std_logic_vector(to_unsigned(165, 8)),
	239 => std_logic_vector(to_unsigned(166, 8)),
	240 => std_logic_vector(to_unsigned(175, 8)),
	241 => std_logic_vector(to_unsigned(164, 8)),
	242 => std_logic_vector(to_unsigned(171, 8)),
	243 => std_logic_vector(to_unsigned(165, 8)),
	244 => std_logic_vector(to_unsigned(173, 8)),
	245 => std_logic_vector(to_unsigned(166, 8)),
	246 => std_logic_vector(to_unsigned(174, 8)),
	247 => std_logic_vector(to_unsigned(172, 8)),
	248 => std_logic_vector(to_unsigned(171, 8)),
	249 => std_logic_vector(to_unsigned(165, 8)),
	250 => std_logic_vector(to_unsigned(171, 8)),
	251 => std_logic_vector(to_unsigned(173, 8)),
	252 => std_logic_vector(to_unsigned(166, 8)),
	253 => std_logic_vector(to_unsigned(172, 8)),
	254 => std_logic_vector(to_unsigned(162, 8)),
	255 => std_logic_vector(to_unsigned(162, 8)),
	256 => std_logic_vector(to_unsigned(168, 8)),
	257 => std_logic_vector(to_unsigned(175, 8)),
	258 => std_logic_vector(to_unsigned(171, 8)),
	259 => std_logic_vector(to_unsigned(169, 8)),
	260 => std_logic_vector(to_unsigned(176, 8)),
	261 => std_logic_vector(to_unsigned(163, 8)),
	262 => std_logic_vector(to_unsigned(168, 8)),
	263 => std_logic_vector(to_unsigned(172, 8)),
	264 => std_logic_vector(to_unsigned(165, 8)),
	265 => std_logic_vector(to_unsigned(175, 8)),
	266 => std_logic_vector(to_unsigned(171, 8)),
	267 => std_logic_vector(to_unsigned(172, 8)),
	268 => std_logic_vector(to_unsigned(172, 8)),
	269 => std_logic_vector(to_unsigned(171, 8)),
	270 => std_logic_vector(to_unsigned(168, 8)),
	271 => std_logic_vector(to_unsigned(173, 8)),
	272 => std_logic_vector(to_unsigned(167, 8)),
	273 => std_logic_vector(to_unsigned(173, 8)),
	274 => std_logic_vector(to_unsigned(166, 8)),
	275 => std_logic_vector(to_unsigned(162, 8)),
	276 => std_logic_vector(to_unsigned(167, 8)),
	277 => std_logic_vector(to_unsigned(175, 8)),
	278 => std_logic_vector(to_unsigned(172, 8)),
	279 => std_logic_vector(to_unsigned(172, 8)),
	280 => std_logic_vector(to_unsigned(169, 8)),
	281 => std_logic_vector(to_unsigned(174, 8)),
	282 => std_logic_vector(to_unsigned(168, 8)),
	283 => std_logic_vector(to_unsigned(169, 8)),
	284 => std_logic_vector(to_unsigned(170, 8)),
	285 => std_logic_vector(to_unsigned(168, 8)),
	286 => std_logic_vector(to_unsigned(176, 8)),
	287 => std_logic_vector(to_unsigned(165, 8)),
	288 => std_logic_vector(to_unsigned(175, 8)),
	289 => std_logic_vector(to_unsigned(171, 8)),
	290 => std_logic_vector(to_unsigned(164, 8)),
	291 => std_logic_vector(to_unsigned(170, 8)),
	292 => std_logic_vector(to_unsigned(168, 8)),
	293 => std_logic_vector(to_unsigned(173, 8)),
	294 => std_logic_vector(to_unsigned(168, 8)),
	295 => std_logic_vector(to_unsigned(174, 8)),
	296 => std_logic_vector(to_unsigned(164, 8)),
	297 => std_logic_vector(to_unsigned(171, 8)),
	298 => std_logic_vector(to_unsigned(169, 8)),
	299 => std_logic_vector(to_unsigned(176, 8)),
	300 => std_logic_vector(to_unsigned(166, 8)),
	301 => std_logic_vector(to_unsigned(168, 8)),
	302 => std_logic_vector(to_unsigned(165, 8)),
	303 => std_logic_vector(to_unsigned(166, 8)),
	304 => std_logic_vector(to_unsigned(162, 8)),
	305 => std_logic_vector(to_unsigned(165, 8)),
	306 => std_logic_vector(to_unsigned(175, 8)),
	307 => std_logic_vector(to_unsigned(163, 8)),
	308 => std_logic_vector(to_unsigned(167, 8)),
	309 => std_logic_vector(to_unsigned(163, 8)),
	310 => std_logic_vector(to_unsigned(172, 8)),
	311 => std_logic_vector(to_unsigned(171, 8)),
	312 => std_logic_vector(to_unsigned(176, 8)),
	313 => std_logic_vector(to_unsigned(165, 8)),
	314 => std_logic_vector(to_unsigned(174, 8)),
	315 => std_logic_vector(to_unsigned(168, 8)),
	316 => std_logic_vector(to_unsigned(167, 8)),
	317 => std_logic_vector(to_unsigned(171, 8)),
	318 => std_logic_vector(to_unsigned(162, 8)),
	319 => std_logic_vector(to_unsigned(165, 8)),
	320 => std_logic_vector(to_unsigned(172, 8)),
	321 => std_logic_vector(to_unsigned(166, 8)),
	322 => std_logic_vector(to_unsigned(162, 8)),
	323 => std_logic_vector(to_unsigned(173, 8)),
	324 => std_logic_vector(to_unsigned(167, 8)),
	325 => std_logic_vector(to_unsigned(167, 8)),
	326 => std_logic_vector(to_unsigned(175, 8)),
	327 => std_logic_vector(to_unsigned(167, 8)),
	328 => std_logic_vector(to_unsigned(176, 8)),
	329 => std_logic_vector(to_unsigned(170, 8)),
	330 => std_logic_vector(to_unsigned(166, 8)),
	331 => std_logic_vector(to_unsigned(162, 8)),
	332 => std_logic_vector(to_unsigned(164, 8)),
	333 => std_logic_vector(to_unsigned(171, 8)),
	334 => std_logic_vector(to_unsigned(164, 8)),
	335 => std_logic_vector(to_unsigned(172, 8)),
	336 => std_logic_vector(to_unsigned(176, 8)),
	337 => std_logic_vector(to_unsigned(169, 8)),
	338 => std_logic_vector(to_unsigned(166, 8)),
	339 => std_logic_vector(to_unsigned(175, 8)),
	340 => std_logic_vector(to_unsigned(168, 8)),
	341 => std_logic_vector(to_unsigned(175, 8)),
	342 => std_logic_vector(to_unsigned(176, 8)),
	343 => std_logic_vector(to_unsigned(173, 8)),
	344 => std_logic_vector(to_unsigned(169, 8)),
	345 => std_logic_vector(to_unsigned(173, 8)),
	346 => std_logic_vector(to_unsigned(162, 8)),
	347 => std_logic_vector(to_unsigned(165, 8)),
	348 => std_logic_vector(to_unsigned(172, 8)),
	349 => std_logic_vector(to_unsigned(172, 8)),
	350 => std_logic_vector(to_unsigned(162, 8)),
	351 => std_logic_vector(to_unsigned(169, 8)),
	352 => std_logic_vector(to_unsigned(165, 8)),
	353 => std_logic_vector(to_unsigned(174, 8)),
	354 => std_logic_vector(to_unsigned(165, 8)),
	355 => std_logic_vector(to_unsigned(162, 8)),
	356 => std_logic_vector(to_unsigned(171, 8)),
	357 => std_logic_vector(to_unsigned(173, 8)),
	358 => std_logic_vector(to_unsigned(172, 8)),
	359 => std_logic_vector(to_unsigned(174, 8)),
	360 => std_logic_vector(to_unsigned(172, 8)),
	361 => std_logic_vector(to_unsigned(170, 8)),
	362 => std_logic_vector(to_unsigned(167, 8)),
	363 => std_logic_vector(to_unsigned(165, 8)),
	364 => std_logic_vector(to_unsigned(170, 8)),
	365 => std_logic_vector(to_unsigned(174, 8)),
	366 => std_logic_vector(to_unsigned(166, 8)),
	367 => std_logic_vector(to_unsigned(166, 8)),
	368 => std_logic_vector(to_unsigned(176, 8)),
	369 => std_logic_vector(to_unsigned(174, 8)),
	370 => std_logic_vector(to_unsigned(175, 8)),
	371 => std_logic_vector(to_unsigned(176, 8)),
	372 => std_logic_vector(to_unsigned(176, 8)),
	373 => std_logic_vector(to_unsigned(174, 8)),
	374 => std_logic_vector(to_unsigned(171, 8)),
	375 => std_logic_vector(to_unsigned(164, 8)),
	376 => std_logic_vector(to_unsigned(167, 8)),
	377 => std_logic_vector(to_unsigned(172, 8)),
	378 => std_logic_vector(to_unsigned(172, 8)),
	379 => std_logic_vector(to_unsigned(171, 8)),
	380 => std_logic_vector(to_unsigned(169, 8)),
	381 => std_logic_vector(to_unsigned(164, 8)),
	382 => std_logic_vector(to_unsigned(163, 8)),
	383 => std_logic_vector(to_unsigned(167, 8)),
	384 => std_logic_vector(to_unsigned(170, 8)),
	385 => std_logic_vector(to_unsigned(170, 8)),
	386 => std_logic_vector(to_unsigned(176, 8)),
	387 => std_logic_vector(to_unsigned(170, 8)),
	388 => std_logic_vector(to_unsigned(169, 8)),
	389 => std_logic_vector(to_unsigned(176, 8)),
	390 => std_logic_vector(to_unsigned(169, 8)),
	391 => std_logic_vector(to_unsigned(171, 8)),
	392 => std_logic_vector(to_unsigned(173, 8)),
	393 => std_logic_vector(to_unsigned(169, 8)),
	394 => std_logic_vector(to_unsigned(173, 8)),
	395 => std_logic_vector(to_unsigned(164, 8)),
	396 => std_logic_vector(to_unsigned(164, 8)),
	397 => std_logic_vector(to_unsigned(176, 8)),
	398 => std_logic_vector(to_unsigned(174, 8)),
	399 => std_logic_vector(to_unsigned(173, 8)),
	400 => std_logic_vector(to_unsigned(164, 8)),
	401 => std_logic_vector(to_unsigned(169, 8)),
	402 => std_logic_vector(to_unsigned(172, 8)),
	403 => std_logic_vector(to_unsigned(168, 8)),
	404 => std_logic_vector(to_unsigned(174, 8)),
	405 => std_logic_vector(to_unsigned(174, 8)),
	406 => std_logic_vector(to_unsigned(163, 8)),
	407 => std_logic_vector(to_unsigned(164, 8)),
	408 => std_logic_vector(to_unsigned(172, 8)),
	409 => std_logic_vector(to_unsigned(165, 8)),
	410 => std_logic_vector(to_unsigned(163, 8)),
	411 => std_logic_vector(to_unsigned(175, 8)),
	412 => std_logic_vector(to_unsigned(175, 8)),
	413 => std_logic_vector(to_unsigned(163, 8)),
	414 => std_logic_vector(to_unsigned(166, 8)),
	415 => std_logic_vector(to_unsigned(163, 8)),
	416 => std_logic_vector(to_unsigned(174, 8)),
	417 => std_logic_vector(to_unsigned(171, 8)),
	418 => std_logic_vector(to_unsigned(165, 8)),
	419 => std_logic_vector(to_unsigned(169, 8)),
	420 => std_logic_vector(to_unsigned(176, 8)),
	421 => std_logic_vector(to_unsigned(162, 8)),
	422 => std_logic_vector(to_unsigned(168, 8)),
	423 => std_logic_vector(to_unsigned(164, 8)),
	424 => std_logic_vector(to_unsigned(169, 8)),
	425 => std_logic_vector(to_unsigned(162, 8)),
	426 => std_logic_vector(to_unsigned(169, 8)),
	427 => std_logic_vector(to_unsigned(175, 8)),
	428 => std_logic_vector(to_unsigned(168, 8)),
	429 => std_logic_vector(to_unsigned(173, 8)),
	430 => std_logic_vector(to_unsigned(169, 8)),
	431 => std_logic_vector(to_unsigned(166, 8)),
	432 => std_logic_vector(to_unsigned(168, 8)),
	433 => std_logic_vector(to_unsigned(172, 8)),
	434 => std_logic_vector(to_unsigned(167, 8)),
	435 => std_logic_vector(to_unsigned(170, 8)),
	436 => std_logic_vector(to_unsigned(168, 8)),
	437 => std_logic_vector(to_unsigned(176, 8)),
	438 => std_logic_vector(to_unsigned(168, 8)),
	439 => std_logic_vector(to_unsigned(173, 8)),
	440 => std_logic_vector(to_unsigned(176, 8)),
	441 => std_logic_vector(to_unsigned(172, 8)),
	442 => std_logic_vector(to_unsigned(164, 8)),
	443 => std_logic_vector(to_unsigned(168, 8)),
	444 => std_logic_vector(to_unsigned(168, 8)),
	445 => std_logic_vector(to_unsigned(163, 8)),
	446 => std_logic_vector(to_unsigned(175, 8)),
	447 => std_logic_vector(to_unsigned(175, 8)),
	448 => std_logic_vector(to_unsigned(175, 8)),
	449 => std_logic_vector(to_unsigned(168, 8)),
	450 => std_logic_vector(to_unsigned(172, 8)),
	451 => std_logic_vector(to_unsigned(162, 8)),
	452 => std_logic_vector(to_unsigned(162, 8)),
	453 => std_logic_vector(to_unsigned(169, 8)),
	454 => std_logic_vector(to_unsigned(176, 8)),
	455 => std_logic_vector(to_unsigned(164, 8)),
	456 => std_logic_vector(to_unsigned(162, 8)),
	457 => std_logic_vector(to_unsigned(169, 8)),
	458 => std_logic_vector(to_unsigned(167, 8)),
	459 => std_logic_vector(to_unsigned(171, 8)),
	460 => std_logic_vector(to_unsigned(169, 8)),
	461 => std_logic_vector(to_unsigned(170, 8)),
	462 => std_logic_vector(to_unsigned(170, 8)),
	463 => std_logic_vector(to_unsigned(174, 8)),
	464 => std_logic_vector(to_unsigned(176, 8)),
	465 => std_logic_vector(to_unsigned(168, 8)),
	466 => std_logic_vector(to_unsigned(166, 8)),
	467 => std_logic_vector(to_unsigned(168, 8)),
	468 => std_logic_vector(to_unsigned(173, 8)),
	469 => std_logic_vector(to_unsigned(170, 8)),
	470 => std_logic_vector(to_unsigned(176, 8)),
	471 => std_logic_vector(to_unsigned(173, 8)),
	472 => std_logic_vector(to_unsigned(165, 8)),
	473 => std_logic_vector(to_unsigned(174, 8)),
	474 => std_logic_vector(to_unsigned(167, 8)),
	475 => std_logic_vector(to_unsigned(172, 8)),
	476 => std_logic_vector(to_unsigned(162, 8)),
	477 => std_logic_vector(to_unsigned(165, 8)),
	478 => std_logic_vector(to_unsigned(162, 8)),
	479 => std_logic_vector(to_unsigned(172, 8)),
	480 => std_logic_vector(to_unsigned(173, 8)),
	481 => std_logic_vector(to_unsigned(164, 8)),
	482 => std_logic_vector(to_unsigned(166, 8)),
	483 => std_logic_vector(to_unsigned(169, 8)),
	484 => std_logic_vector(to_unsigned(170, 8)),
	485 => std_logic_vector(to_unsigned(171, 8)),
	486 => std_logic_vector(to_unsigned(169, 8)),
	487 => std_logic_vector(to_unsigned(173, 8)),
	488 => std_logic_vector(to_unsigned(162, 8)),
	489 => std_logic_vector(to_unsigned(167, 8)),
	490 => std_logic_vector(to_unsigned(175, 8)),
	491 => std_logic_vector(to_unsigned(167, 8)),
	492 => std_logic_vector(to_unsigned(166, 8)),
	493 => std_logic_vector(to_unsigned(174, 8)),
	494 => std_logic_vector(to_unsigned(173, 8)),
	495 => std_logic_vector(to_unsigned(174, 8)),
	496 => std_logic_vector(to_unsigned(164, 8)),
	497 => std_logic_vector(to_unsigned(172, 8)),
	498 => std_logic_vector(to_unsigned(166, 8)),
	499 => std_logic_vector(to_unsigned(176, 8)),
	500 => std_logic_vector(to_unsigned(173, 8)),
	501 => std_logic_vector(to_unsigned(163, 8)),
	502 => std_logic_vector(to_unsigned(172, 8)),
	503 => std_logic_vector(to_unsigned(170, 8)),
	504 => std_logic_vector(to_unsigned(163, 8)),
	505 => std_logic_vector(to_unsigned(174, 8)),
	506 => std_logic_vector(to_unsigned(173, 8)),
	507 => std_logic_vector(to_unsigned(167, 8)),
	508 => std_logic_vector(to_unsigned(176, 8)),
	509 => std_logic_vector(to_unsigned(164, 8)),
	510 => std_logic_vector(to_unsigned(165, 8)),
	511 => std_logic_vector(to_unsigned(175, 8)),
	512 => std_logic_vector(to_unsigned(162, 8)),
	513 => std_logic_vector(to_unsigned(166, 8)),
	514 => std_logic_vector(to_unsigned(174, 8)),
	515 => std_logic_vector(to_unsigned(168, 8)),
	516 => std_logic_vector(to_unsigned(171, 8)),
	517 => std_logic_vector(to_unsigned(170, 8)),
	518 => std_logic_vector(to_unsigned(174, 8)),
	519 => std_logic_vector(to_unsigned(170, 8)),
	520 => std_logic_vector(to_unsigned(165, 8)),
	521 => std_logic_vector(to_unsigned(164, 8)),
	522 => std_logic_vector(to_unsigned(174, 8)),
	523 => std_logic_vector(to_unsigned(165, 8)),
	524 => std_logic_vector(to_unsigned(171, 8)),
	525 => std_logic_vector(to_unsigned(175, 8)),
	526 => std_logic_vector(to_unsigned(175, 8)),
	527 => std_logic_vector(to_unsigned(162, 8)),
	528 => std_logic_vector(to_unsigned(172, 8)),
	529 => std_logic_vector(to_unsigned(166, 8)),
	530 => std_logic_vector(to_unsigned(163, 8)),
	531 => std_logic_vector(to_unsigned(176, 8)),
	532 => std_logic_vector(to_unsigned(165, 8)),
	533 => std_logic_vector(to_unsigned(166, 8)),
	534 => std_logic_vector(to_unsigned(165, 8)),
	535 => std_logic_vector(to_unsigned(169, 8)),
	536 => std_logic_vector(to_unsigned(174, 8)),
	537 => std_logic_vector(to_unsigned(165, 8)),
	538 => std_logic_vector(to_unsigned(165, 8)),
	539 => std_logic_vector(to_unsigned(162, 8)),
	540 => std_logic_vector(to_unsigned(170, 8)),
	541 => std_logic_vector(to_unsigned(174, 8)),
	542 => std_logic_vector(to_unsigned(163, 8)),
	543 => std_logic_vector(to_unsigned(174, 8)),
	544 => std_logic_vector(to_unsigned(176, 8)),
	545 => std_logic_vector(to_unsigned(168, 8)),
	546 => std_logic_vector(to_unsigned(171, 8)),
	547 => std_logic_vector(to_unsigned(176, 8)),
	548 => std_logic_vector(to_unsigned(167, 8)),
	549 => std_logic_vector(to_unsigned(163, 8)),
	550 => std_logic_vector(to_unsigned(170, 8)),
	551 => std_logic_vector(to_unsigned(170, 8)),
	552 => std_logic_vector(to_unsigned(163, 8)),
	553 => std_logic_vector(to_unsigned(167, 8)),
	554 => std_logic_vector(to_unsigned(171, 8)),
	555 => std_logic_vector(to_unsigned(175, 8)),
	556 => std_logic_vector(to_unsigned(169, 8)),
	557 => std_logic_vector(to_unsigned(175, 8)),
	558 => std_logic_vector(to_unsigned(168, 8)),
	559 => std_logic_vector(to_unsigned(173, 8)),
	560 => std_logic_vector(to_unsigned(176, 8)),
	561 => std_logic_vector(to_unsigned(162, 8)),
	562 => std_logic_vector(to_unsigned(172, 8)),
	563 => std_logic_vector(to_unsigned(174, 8)),
	564 => std_logic_vector(to_unsigned(169, 8)),
	565 => std_logic_vector(to_unsigned(174, 8)),
	566 => std_logic_vector(to_unsigned(175, 8)),
	567 => std_logic_vector(to_unsigned(170, 8)),
	568 => std_logic_vector(to_unsigned(174, 8)),
	569 => std_logic_vector(to_unsigned(172, 8)),
	570 => std_logic_vector(to_unsigned(169, 8)),
	571 => std_logic_vector(to_unsigned(174, 8)),
	572 => std_logic_vector(to_unsigned(173, 8)),
	573 => std_logic_vector(to_unsigned(172, 8)),
	574 => std_logic_vector(to_unsigned(174, 8)),
	575 => std_logic_vector(to_unsigned(164, 8)),
	576 => std_logic_vector(to_unsigned(167, 8)),
	577 => std_logic_vector(to_unsigned(169, 8)),
	578 => std_logic_vector(to_unsigned(164, 8)),
	579 => std_logic_vector(to_unsigned(166, 8)),
	580 => std_logic_vector(to_unsigned(162, 8)),
	581 => std_logic_vector(to_unsigned(163, 8)),
	582 => std_logic_vector(to_unsigned(163, 8)),
	583 => std_logic_vector(to_unsigned(171, 8)),
	584 => std_logic_vector(to_unsigned(169, 8)),
	585 => std_logic_vector(to_unsigned(171, 8)),
	586 => std_logic_vector(to_unsigned(165, 8)),
	587 => std_logic_vector(to_unsigned(172, 8)),
	588 => std_logic_vector(to_unsigned(163, 8)),
	589 => std_logic_vector(to_unsigned(164, 8)),
	590 => std_logic_vector(to_unsigned(164, 8)),
	591 => std_logic_vector(to_unsigned(166, 8)),
	592 => std_logic_vector(to_unsigned(169, 8)),
	593 => std_logic_vector(to_unsigned(170, 8)),
	594 => std_logic_vector(to_unsigned(168, 8)),
	595 => std_logic_vector(to_unsigned(167, 8)),
	596 => std_logic_vector(to_unsigned(162, 8)),
	597 => std_logic_vector(to_unsigned(162, 8)),
	598 => std_logic_vector(to_unsigned(174, 8)),
	599 => std_logic_vector(to_unsigned(169, 8)),
	600 => std_logic_vector(to_unsigned(162, 8)),
	601 => std_logic_vector(to_unsigned(164, 8)),
	602 => std_logic_vector(to_unsigned(175, 8)),
	603 => std_logic_vector(to_unsigned(166, 8)),
	604 => std_logic_vector(to_unsigned(164, 8)),
	605 => std_logic_vector(to_unsigned(164, 8)),
	606 => std_logic_vector(to_unsigned(173, 8)),
	607 => std_logic_vector(to_unsigned(163, 8)),
	608 => std_logic_vector(to_unsigned(174, 8)),
	609 => std_logic_vector(to_unsigned(164, 8)),
	610 => std_logic_vector(to_unsigned(165, 8)),
	611 => std_logic_vector(to_unsigned(175, 8)),
	612 => std_logic_vector(to_unsigned(174, 8)),
	613 => std_logic_vector(to_unsigned(166, 8)),
	614 => std_logic_vector(to_unsigned(166, 8)),
	615 => std_logic_vector(to_unsigned(172, 8)),
	616 => std_logic_vector(to_unsigned(162, 8)),
	617 => std_logic_vector(to_unsigned(165, 8)),
	618 => std_logic_vector(to_unsigned(174, 8)),
	619 => std_logic_vector(to_unsigned(174, 8)),
	620 => std_logic_vector(to_unsigned(174, 8)),
	621 => std_logic_vector(to_unsigned(176, 8)),
	622 => std_logic_vector(to_unsigned(173, 8)),
	623 => std_logic_vector(to_unsigned(163, 8)),
	624 => std_logic_vector(to_unsigned(168, 8)),
	625 => std_logic_vector(to_unsigned(173, 8)),
	626 => std_logic_vector(to_unsigned(168, 8)),
	627 => std_logic_vector(to_unsigned(167, 8)),
	628 => std_logic_vector(to_unsigned(171, 8)),
	629 => std_logic_vector(to_unsigned(165, 8)),
	630 => std_logic_vector(to_unsigned(166, 8)),
	631 => std_logic_vector(to_unsigned(171, 8)),
	632 => std_logic_vector(to_unsigned(170, 8)),
	633 => std_logic_vector(to_unsigned(166, 8)),
	634 => std_logic_vector(to_unsigned(176, 8)),
	635 => std_logic_vector(to_unsigned(170, 8)),
	636 => std_logic_vector(to_unsigned(175, 8)),
	637 => std_logic_vector(to_unsigned(163, 8)),
	638 => std_logic_vector(to_unsigned(167, 8)),
	639 => std_logic_vector(to_unsigned(169, 8)),
	640 => std_logic_vector(to_unsigned(168, 8)),
	641 => std_logic_vector(to_unsigned(165, 8)),
	642 => std_logic_vector(to_unsigned(176, 8)),
	643 => std_logic_vector(to_unsigned(175, 8)),
	644 => std_logic_vector(to_unsigned(176, 8)),
	645 => std_logic_vector(to_unsigned(165, 8)),
	646 => std_logic_vector(to_unsigned(175, 8)),
	647 => std_logic_vector(to_unsigned(168, 8)),
	648 => std_logic_vector(to_unsigned(167, 8)),
	649 => std_logic_vector(to_unsigned(172, 8)),
	650 => std_logic_vector(to_unsigned(162, 8)),
	651 => std_logic_vector(to_unsigned(174, 8)),
	652 => std_logic_vector(to_unsigned(175, 8)),
	653 => std_logic_vector(to_unsigned(174, 8)),
	654 => std_logic_vector(to_unsigned(170, 8)),
	655 => std_logic_vector(to_unsigned(164, 8)),
	656 => std_logic_vector(to_unsigned(167, 8)),
	657 => std_logic_vector(to_unsigned(162, 8)),
	658 => std_logic_vector(to_unsigned(162, 8)),
	659 => std_logic_vector(to_unsigned(170, 8)),
	660 => std_logic_vector(to_unsigned(171, 8)),
	661 => std_logic_vector(to_unsigned(169, 8)),
	662 => std_logic_vector(to_unsigned(175, 8)),
	663 => std_logic_vector(to_unsigned(168, 8)),
	664 => std_logic_vector(to_unsigned(169, 8)),
	665 => std_logic_vector(to_unsigned(167, 8)),
	666 => std_logic_vector(to_unsigned(171, 8)),
	667 => std_logic_vector(to_unsigned(173, 8)),
	668 => std_logic_vector(to_unsigned(174, 8)),
	669 => std_logic_vector(to_unsigned(172, 8)),
	670 => std_logic_vector(to_unsigned(167, 8)),
	671 => std_logic_vector(to_unsigned(173, 8)),
	672 => std_logic_vector(to_unsigned(167, 8)),
	673 => std_logic_vector(to_unsigned(174, 8)),
	674 => std_logic_vector(to_unsigned(164, 8)),
	675 => std_logic_vector(to_unsigned(166, 8)),
	676 => std_logic_vector(to_unsigned(169, 8)),
	677 => std_logic_vector(to_unsigned(165, 8)),
	678 => std_logic_vector(to_unsigned(162, 8)),
	679 => std_logic_vector(to_unsigned(170, 8)),
	680 => std_logic_vector(to_unsigned(164, 8)),
	681 => std_logic_vector(to_unsigned(169, 8)),
	682 => std_logic_vector(to_unsigned(163, 8)),
	683 => std_logic_vector(to_unsigned(166, 8)),
	684 => std_logic_vector(to_unsigned(163, 8)),
	685 => std_logic_vector(to_unsigned(172, 8)),
	686 => std_logic_vector(to_unsigned(164, 8)),
	687 => std_logic_vector(to_unsigned(171, 8)),
	688 => std_logic_vector(to_unsigned(174, 8)),
	689 => std_logic_vector(to_unsigned(173, 8)),
	690 => std_logic_vector(to_unsigned(165, 8)),
	691 => std_logic_vector(to_unsigned(167, 8)),
	692 => std_logic_vector(to_unsigned(162, 8)),
	693 => std_logic_vector(to_unsigned(176, 8)),
	694 => std_logic_vector(to_unsigned(162, 8)),
	695 => std_logic_vector(to_unsigned(163, 8)),
	696 => std_logic_vector(to_unsigned(171, 8)),
	697 => std_logic_vector(to_unsigned(175, 8)),
	698 => std_logic_vector(to_unsigned(171, 8)),
	699 => std_logic_vector(to_unsigned(175, 8)),
	700 => std_logic_vector(to_unsigned(167, 8)),
	701 => std_logic_vector(to_unsigned(167, 8)),
	702 => std_logic_vector(to_unsigned(162, 8)),
	703 => std_logic_vector(to_unsigned(171, 8)),
	704 => std_logic_vector(to_unsigned(173, 8)),
	705 => std_logic_vector(to_unsigned(170, 8)),
	706 => std_logic_vector(to_unsigned(168, 8)),
	707 => std_logic_vector(to_unsigned(170, 8)),
	708 => std_logic_vector(to_unsigned(163, 8)),
	709 => std_logic_vector(to_unsigned(164, 8)),
	710 => std_logic_vector(to_unsigned(173, 8)),
	711 => std_logic_vector(to_unsigned(171, 8)),
	712 => std_logic_vector(to_unsigned(170, 8)),
	713 => std_logic_vector(to_unsigned(168, 8)),
	714 => std_logic_vector(to_unsigned(172, 8)),
	715 => std_logic_vector(to_unsigned(162, 8)),
	716 => std_logic_vector(to_unsigned(176, 8)),
	717 => std_logic_vector(to_unsigned(164, 8)),
	718 => std_logic_vector(to_unsigned(175, 8)),
	719 => std_logic_vector(to_unsigned(163, 8)),
	720 => std_logic_vector(to_unsigned(173, 8)),
	721 => std_logic_vector(to_unsigned(168, 8)),
	722 => std_logic_vector(to_unsigned(168, 8)),
	723 => std_logic_vector(to_unsigned(175, 8)),
	724 => std_logic_vector(to_unsigned(172, 8)),
	725 => std_logic_vector(to_unsigned(169, 8)),
	726 => std_logic_vector(to_unsigned(169, 8)),
	727 => std_logic_vector(to_unsigned(166, 8)),
	728 => std_logic_vector(to_unsigned(173, 8)),
	729 => std_logic_vector(to_unsigned(175, 8)),
	730 => std_logic_vector(to_unsigned(170, 8)),
	731 => std_logic_vector(to_unsigned(172, 8)),
	732 => std_logic_vector(to_unsigned(168, 8)),
	733 => std_logic_vector(to_unsigned(168, 8)),
	734 => std_logic_vector(to_unsigned(170, 8)),
	735 => std_logic_vector(to_unsigned(175, 8)),
	736 => std_logic_vector(to_unsigned(163, 8)),
	737 => std_logic_vector(to_unsigned(167, 8)),
	738 => std_logic_vector(to_unsigned(164, 8)),
	739 => std_logic_vector(to_unsigned(170, 8)),
	740 => std_logic_vector(to_unsigned(165, 8)),
	741 => std_logic_vector(to_unsigned(165, 8)),
	742 => std_logic_vector(to_unsigned(167, 8)),
	743 => std_logic_vector(to_unsigned(165, 8)),
	744 => std_logic_vector(to_unsigned(162, 8)),
	745 => std_logic_vector(to_unsigned(162, 8)),
	746 => std_logic_vector(to_unsigned(164, 8)),
	747 => std_logic_vector(to_unsigned(168, 8)),
	748 => std_logic_vector(to_unsigned(166, 8)),
	749 => std_logic_vector(to_unsigned(163, 8)),
	750 => std_logic_vector(to_unsigned(162, 8)),
	751 => std_logic_vector(to_unsigned(164, 8)),
	752 => std_logic_vector(to_unsigned(167, 8)),
	753 => std_logic_vector(to_unsigned(167, 8)),
	754 => std_logic_vector(to_unsigned(176, 8)),
	755 => std_logic_vector(to_unsigned(170, 8)),
	756 => std_logic_vector(to_unsigned(164, 8)),
	757 => std_logic_vector(to_unsigned(167, 8)),
	758 => std_logic_vector(to_unsigned(173, 8)),
	759 => std_logic_vector(to_unsigned(174, 8)),
	760 => std_logic_vector(to_unsigned(173, 8)),
	761 => std_logic_vector(to_unsigned(167, 8)),
	762 => std_logic_vector(to_unsigned(172, 8)),
	763 => std_logic_vector(to_unsigned(171, 8)),
	764 => std_logic_vector(to_unsigned(169, 8)),
	765 => std_logic_vector(to_unsigned(166, 8)),
	766 => std_logic_vector(to_unsigned(168, 8)),
	767 => std_logic_vector(to_unsigned(162, 8)),
	768 => std_logic_vector(to_unsigned(167, 8)),
	769 => std_logic_vector(to_unsigned(165, 8)),
	770 => std_logic_vector(to_unsigned(163, 8)),
	771 => std_logic_vector(to_unsigned(172, 8)),
	772 => std_logic_vector(to_unsigned(167, 8)),
	773 => std_logic_vector(to_unsigned(176, 8)),
	774 => std_logic_vector(to_unsigned(175, 8)),
	775 => std_logic_vector(to_unsigned(163, 8)),
	776 => std_logic_vector(to_unsigned(165, 8)),
	777 => std_logic_vector(to_unsigned(164, 8)),
	778 => std_logic_vector(to_unsigned(163, 8)),
	779 => std_logic_vector(to_unsigned(171, 8)),
	780 => std_logic_vector(to_unsigned(171, 8)),
	781 => std_logic_vector(to_unsigned(173, 8)),
	782 => std_logic_vector(to_unsigned(166, 8)),
	783 => std_logic_vector(to_unsigned(174, 8)),
	784 => std_logic_vector(to_unsigned(170, 8)),
	785 => std_logic_vector(to_unsigned(172, 8)),
	786 => std_logic_vector(to_unsigned(172, 8)),
	787 => std_logic_vector(to_unsigned(171, 8)),
	788 => std_logic_vector(to_unsigned(168, 8)),
	789 => std_logic_vector(to_unsigned(169, 8)),
	790 => std_logic_vector(to_unsigned(173, 8)),
	791 => std_logic_vector(to_unsigned(173, 8)),
	792 => std_logic_vector(to_unsigned(163, 8)),
	793 => std_logic_vector(to_unsigned(174, 8)),
	794 => std_logic_vector(to_unsigned(172, 8)),
	795 => std_logic_vector(to_unsigned(169, 8)),
	796 => std_logic_vector(to_unsigned(162, 8)),
	797 => std_logic_vector(to_unsigned(173, 8)),
	798 => std_logic_vector(to_unsigned(175, 8)),
	799 => std_logic_vector(to_unsigned(168, 8)),
	800 => std_logic_vector(to_unsigned(166, 8)),
	801 => std_logic_vector(to_unsigned(176, 8)),
	802 => std_logic_vector(to_unsigned(176, 8)),
	803 => std_logic_vector(to_unsigned(168, 8)),
	804 => std_logic_vector(to_unsigned(171, 8)),
	805 => std_logic_vector(to_unsigned(174, 8)),
	806 => std_logic_vector(to_unsigned(175, 8)),
	807 => std_logic_vector(to_unsigned(171, 8)),
	808 => std_logic_vector(to_unsigned(170, 8)),
	809 => std_logic_vector(to_unsigned(165, 8)),
	810 => std_logic_vector(to_unsigned(167, 8)),
	811 => std_logic_vector(to_unsigned(170, 8)),
	812 => std_logic_vector(to_unsigned(167, 8)),
	813 => std_logic_vector(to_unsigned(163, 8)),
	814 => std_logic_vector(to_unsigned(165, 8)),
	815 => std_logic_vector(to_unsigned(165, 8)),
	816 => std_logic_vector(to_unsigned(175, 8)),
	817 => std_logic_vector(to_unsigned(169, 8)),
	818 => std_logic_vector(to_unsigned(172, 8)),
	819 => std_logic_vector(to_unsigned(168, 8)),
	820 => std_logic_vector(to_unsigned(165, 8)),
	821 => std_logic_vector(to_unsigned(168, 8)),
	822 => std_logic_vector(to_unsigned(173, 8)),
	823 => std_logic_vector(to_unsigned(162, 8)),
	824 => std_logic_vector(to_unsigned(170, 8)),
	825 => std_logic_vector(to_unsigned(173, 8)),
	826 => std_logic_vector(to_unsigned(162, 8)),
	827 => std_logic_vector(to_unsigned(175, 8)),
	828 => std_logic_vector(to_unsigned(166, 8)),
	829 => std_logic_vector(to_unsigned(173, 8)),
	830 => std_logic_vector(to_unsigned(162, 8)),
	831 => std_logic_vector(to_unsigned(169, 8)),
	832 => std_logic_vector(to_unsigned(163, 8)),
	833 => std_logic_vector(to_unsigned(162, 8)),
	834 => std_logic_vector(to_unsigned(163, 8)),
	835 => std_logic_vector(to_unsigned(172, 8)),
	836 => std_logic_vector(to_unsigned(166, 8)),
	837 => std_logic_vector(to_unsigned(176, 8)),
	838 => std_logic_vector(to_unsigned(171, 8)),
	839 => std_logic_vector(to_unsigned(163, 8)),
	840 => std_logic_vector(to_unsigned(164, 8)),
	841 => std_logic_vector(to_unsigned(176, 8)),
	842 => std_logic_vector(to_unsigned(170, 8)),
	843 => std_logic_vector(to_unsigned(173, 8)),
	844 => std_logic_vector(to_unsigned(167, 8)),
	845 => std_logic_vector(to_unsigned(162, 8)),
	846 => std_logic_vector(to_unsigned(171, 8)),
	847 => std_logic_vector(to_unsigned(165, 8)),
	848 => std_logic_vector(to_unsigned(163, 8)),
	849 => std_logic_vector(to_unsigned(162, 8)),
	850 => std_logic_vector(to_unsigned(168, 8)),
	851 => std_logic_vector(to_unsigned(176, 8)),
	852 => std_logic_vector(to_unsigned(169, 8)),
	853 => std_logic_vector(to_unsigned(174, 8)),
	854 => std_logic_vector(to_unsigned(173, 8)),
	855 => std_logic_vector(to_unsigned(164, 8)),
	856 => std_logic_vector(to_unsigned(172, 8)),
	857 => std_logic_vector(to_unsigned(167, 8)),
	858 => std_logic_vector(to_unsigned(163, 8)),
	859 => std_logic_vector(to_unsigned(169, 8)),
	860 => std_logic_vector(to_unsigned(171, 8)),
	861 => std_logic_vector(to_unsigned(171, 8)),
	862 => std_logic_vector(to_unsigned(163, 8)),
	863 => std_logic_vector(to_unsigned(171, 8)),
	864 => std_logic_vector(to_unsigned(166, 8)),
	865 => std_logic_vector(to_unsigned(175, 8)),
	866 => std_logic_vector(to_unsigned(174, 8)),
	867 => std_logic_vector(to_unsigned(176, 8)),
	868 => std_logic_vector(to_unsigned(170, 8)),
	869 => std_logic_vector(to_unsigned(168, 8)),
	870 => std_logic_vector(to_unsigned(176, 8)),
	871 => std_logic_vector(to_unsigned(166, 8)),
	872 => std_logic_vector(to_unsigned(162, 8)),
	873 => std_logic_vector(to_unsigned(170, 8)),
	874 => std_logic_vector(to_unsigned(163, 8)),
	875 => std_logic_vector(to_unsigned(163, 8)),
	876 => std_logic_vector(to_unsigned(166, 8)),
	877 => std_logic_vector(to_unsigned(173, 8)),
	878 => std_logic_vector(to_unsigned(170, 8)),
	879 => std_logic_vector(to_unsigned(162, 8)),
	880 => std_logic_vector(to_unsigned(164, 8)),
	881 => std_logic_vector(to_unsigned(172, 8)),
	882 => std_logic_vector(to_unsigned(165, 8)),
	883 => std_logic_vector(to_unsigned(175, 8)),
	884 => std_logic_vector(to_unsigned(165, 8)),
	885 => std_logic_vector(to_unsigned(175, 8)),
	886 => std_logic_vector(to_unsigned(162, 8)),
	887 => std_logic_vector(to_unsigned(171, 8)),
	888 => std_logic_vector(to_unsigned(166, 8)),
	889 => std_logic_vector(to_unsigned(163, 8)),
	890 => std_logic_vector(to_unsigned(169, 8)),
	891 => std_logic_vector(to_unsigned(168, 8)),
	892 => std_logic_vector(to_unsigned(167, 8)),
	893 => std_logic_vector(to_unsigned(172, 8)),
	894 => std_logic_vector(to_unsigned(163, 8)),
	895 => std_logic_vector(to_unsigned(175, 8)),
	896 => std_logic_vector(to_unsigned(164, 8)),
	897 => std_logic_vector(to_unsigned(176, 8)),
	898 => std_logic_vector(to_unsigned(162, 8)),
	899 => std_logic_vector(to_unsigned(169, 8)),
	900 => std_logic_vector(to_unsigned(170, 8)),
	901 => std_logic_vector(to_unsigned(164, 8)),
	902 => std_logic_vector(to_unsigned(168, 8)),
	903 => std_logic_vector(to_unsigned(165, 8)),
	904 => std_logic_vector(to_unsigned(167, 8)),
	905 => std_logic_vector(to_unsigned(162, 8)),
	906 => std_logic_vector(to_unsigned(176, 8)),
	907 => std_logic_vector(to_unsigned(163, 8)),
	908 => std_logic_vector(to_unsigned(162, 8)),
	909 => std_logic_vector(to_unsigned(171, 8)),
	910 => std_logic_vector(to_unsigned(169, 8)),
	911 => std_logic_vector(to_unsigned(168, 8)),
	912 => std_logic_vector(to_unsigned(174, 8)),
	913 => std_logic_vector(to_unsigned(174, 8)),
	914 => std_logic_vector(to_unsigned(173, 8)),
	915 => std_logic_vector(to_unsigned(168, 8)),
	916 => std_logic_vector(to_unsigned(166, 8)),
	917 => std_logic_vector(to_unsigned(176, 8)),
	918 => std_logic_vector(to_unsigned(168, 8)),
	919 => std_logic_vector(to_unsigned(165, 8)),
	920 => std_logic_vector(to_unsigned(168, 8)),
	921 => std_logic_vector(to_unsigned(170, 8)),
	922 => std_logic_vector(to_unsigned(176, 8)),
	923 => std_logic_vector(to_unsigned(166, 8)),
	924 => std_logic_vector(to_unsigned(162, 8)),
	925 => std_logic_vector(to_unsigned(166, 8)),
	926 => std_logic_vector(to_unsigned(176, 8)),
	927 => std_logic_vector(to_unsigned(162, 8)),
	928 => std_logic_vector(to_unsigned(163, 8)),
	929 => std_logic_vector(to_unsigned(164, 8)),
	930 => std_logic_vector(to_unsigned(164, 8)),
	931 => std_logic_vector(to_unsigned(163, 8)),
	932 => std_logic_vector(to_unsigned(162, 8)),
	933 => std_logic_vector(to_unsigned(172, 8)),
	934 => std_logic_vector(to_unsigned(164, 8)),
	935 => std_logic_vector(to_unsigned(164, 8)),
	936 => std_logic_vector(to_unsigned(166, 8)),
	937 => std_logic_vector(to_unsigned(169, 8)),
	938 => std_logic_vector(to_unsigned(173, 8)),
	939 => std_logic_vector(to_unsigned(162, 8)),
	940 => std_logic_vector(to_unsigned(168, 8)),
	941 => std_logic_vector(to_unsigned(172, 8)),
	942 => std_logic_vector(to_unsigned(167, 8)),
	943 => std_logic_vector(to_unsigned(171, 8)),
	944 => std_logic_vector(to_unsigned(164, 8)),
	945 => std_logic_vector(to_unsigned(172, 8)),
	946 => std_logic_vector(to_unsigned(169, 8)),
	947 => std_logic_vector(to_unsigned(166, 8)),
	948 => std_logic_vector(to_unsigned(176, 8)),
	949 => std_logic_vector(to_unsigned(167, 8)),
	950 => std_logic_vector(to_unsigned(164, 8)),
	951 => std_logic_vector(to_unsigned(164, 8)),
	952 => std_logic_vector(to_unsigned(172, 8)),
	953 => std_logic_vector(to_unsigned(162, 8)),
	954 => std_logic_vector(to_unsigned(167, 8)),
	955 => std_logic_vector(to_unsigned(162, 8)),
	956 => std_logic_vector(to_unsigned(164, 8)),
	957 => std_logic_vector(to_unsigned(174, 8)),
	958 => std_logic_vector(to_unsigned(167, 8)),
	959 => std_logic_vector(to_unsigned(171, 8)),
	960 => std_logic_vector(to_unsigned(168, 8)),
	961 => std_logic_vector(to_unsigned(162, 8)),
	962 => std_logic_vector(to_unsigned(167, 8)),
	963 => std_logic_vector(to_unsigned(164, 8)),
	964 => std_logic_vector(to_unsigned(175, 8)),
	965 => std_logic_vector(to_unsigned(176, 8)),
	966 => std_logic_vector(to_unsigned(172, 8)),
	967 => std_logic_vector(to_unsigned(163, 8)),
	968 => std_logic_vector(to_unsigned(168, 8)),
	969 => std_logic_vector(to_unsigned(166, 8)),
	970 => std_logic_vector(to_unsigned(169, 8)),
	971 => std_logic_vector(to_unsigned(165, 8)),
	972 => std_logic_vector(to_unsigned(168, 8)),
	973 => std_logic_vector(to_unsigned(165, 8)),
	974 => std_logic_vector(to_unsigned(163, 8)),
	975 => std_logic_vector(to_unsigned(169, 8)),
	976 => std_logic_vector(to_unsigned(163, 8)),
	977 => std_logic_vector(to_unsigned(169, 8)),
	978 => std_logic_vector(to_unsigned(162, 8)),
	979 => std_logic_vector(to_unsigned(172, 8)),
	980 => std_logic_vector(to_unsigned(168, 8)),
	981 => std_logic_vector(to_unsigned(164, 8)),
	982 => std_logic_vector(to_unsigned(169, 8)),
	983 => std_logic_vector(to_unsigned(171, 8)),
	984 => std_logic_vector(to_unsigned(175, 8)),
	985 => std_logic_vector(to_unsigned(167, 8)),
	986 => std_logic_vector(to_unsigned(165, 8)),
	987 => std_logic_vector(to_unsigned(162, 8)),
	988 => std_logic_vector(to_unsigned(173, 8)),
	989 => std_logic_vector(to_unsigned(175, 8)),
	990 => std_logic_vector(to_unsigned(166, 8)),
	991 => std_logic_vector(to_unsigned(175, 8)),
	992 => std_logic_vector(to_unsigned(165, 8)),
	993 => std_logic_vector(to_unsigned(170, 8)),
	994 => std_logic_vector(to_unsigned(166, 8)),
	995 => std_logic_vector(to_unsigned(168, 8)),
	996 => std_logic_vector(to_unsigned(176, 8)),
	997 => std_logic_vector(to_unsigned(173, 8)),
	998 => std_logic_vector(to_unsigned(173, 8)),
	999 => std_logic_vector(to_unsigned(171, 8)),
	1000 => std_logic_vector(to_unsigned(163, 8)),
	1001 => std_logic_vector(to_unsigned(170, 8)),
	1002 => std_logic_vector(to_unsigned(165, 8)),
	1003 => std_logic_vector(to_unsigned(163, 8)),
	1004 => std_logic_vector(to_unsigned(164, 8)),
	1005 => std_logic_vector(to_unsigned(165, 8)),
	1006 => std_logic_vector(to_unsigned(173, 8)),
	1007 => std_logic_vector(to_unsigned(167, 8)),
	1008 => std_logic_vector(to_unsigned(162, 8)),
	1009 => std_logic_vector(to_unsigned(164, 8)),
	1010 => std_logic_vector(to_unsigned(164, 8)),
	1011 => std_logic_vector(to_unsigned(164, 8)),
	1012 => std_logic_vector(to_unsigned(163, 8)),
	1013 => std_logic_vector(to_unsigned(166, 8)),
	1014 => std_logic_vector(to_unsigned(173, 8)),
	1015 => std_logic_vector(to_unsigned(169, 8)),
	1016 => std_logic_vector(to_unsigned(169, 8)),
	1017 => std_logic_vector(to_unsigned(163, 8)),
	1018 => std_logic_vector(to_unsigned(171, 8)),
	1019 => std_logic_vector(to_unsigned(175, 8)),
	1020 => std_logic_vector(to_unsigned(173, 8)),
	1021 => std_logic_vector(to_unsigned(166, 8)),
	1022 => std_logic_vector(to_unsigned(163, 8)),
	1023 => std_logic_vector(to_unsigned(165, 8)),
	1024 => std_logic_vector(to_unsigned(172, 8)),
	1025 => std_logic_vector(to_unsigned(165, 8)),
	1026 => std_logic_vector(to_unsigned(171, 8)),
	1027 => std_logic_vector(to_unsigned(167, 8)),
	1028 => std_logic_vector(to_unsigned(165, 8)),
	1029 => std_logic_vector(to_unsigned(167, 8)),
	1030 => std_logic_vector(to_unsigned(162, 8)),
	1031 => std_logic_vector(to_unsigned(165, 8)),
	1032 => std_logic_vector(to_unsigned(163, 8)),
	1033 => std_logic_vector(to_unsigned(166, 8)),
	1034 => std_logic_vector(to_unsigned(172, 8)),
	1035 => std_logic_vector(to_unsigned(172, 8)),
	1036 => std_logic_vector(to_unsigned(169, 8)),
	1037 => std_logic_vector(to_unsigned(168, 8)),
	1038 => std_logic_vector(to_unsigned(172, 8)),
	1039 => std_logic_vector(to_unsigned(171, 8)),
	1040 => std_logic_vector(to_unsigned(162, 8)),
	1041 => std_logic_vector(to_unsigned(171, 8)),
	1042 => std_logic_vector(to_unsigned(167, 8)),
	1043 => std_logic_vector(to_unsigned(167, 8)),
	1044 => std_logic_vector(to_unsigned(164, 8)),
	1045 => std_logic_vector(to_unsigned(170, 8)),
	1046 => std_logic_vector(to_unsigned(172, 8)),
	1047 => std_logic_vector(to_unsigned(167, 8)),
	1048 => std_logic_vector(to_unsigned(168, 8)),
	1049 => std_logic_vector(to_unsigned(174, 8)),
	1050 => std_logic_vector(to_unsigned(169, 8)),
	1051 => std_logic_vector(to_unsigned(174, 8)),
	1052 => std_logic_vector(to_unsigned(165, 8)),
	1053 => std_logic_vector(to_unsigned(173, 8)),
	1054 => std_logic_vector(to_unsigned(171, 8)),
	1055 => std_logic_vector(to_unsigned(167, 8)),
	1056 => std_logic_vector(to_unsigned(175, 8)),
	1057 => std_logic_vector(to_unsigned(164, 8)),
	1058 => std_logic_vector(to_unsigned(175, 8)),
	1059 => std_logic_vector(to_unsigned(173, 8)),
	1060 => std_logic_vector(to_unsigned(165, 8)),
	1061 => std_logic_vector(to_unsigned(170, 8)),
	1062 => std_logic_vector(to_unsigned(170, 8)),
	1063 => std_logic_vector(to_unsigned(170, 8)),
	1064 => std_logic_vector(to_unsigned(172, 8)),
	1065 => std_logic_vector(to_unsigned(164, 8)),
	1066 => std_logic_vector(to_unsigned(170, 8)),
	1067 => std_logic_vector(to_unsigned(163, 8)),
	1068 => std_logic_vector(to_unsigned(163, 8)),
	1069 => std_logic_vector(to_unsigned(173, 8)),
	1070 => std_logic_vector(to_unsigned(172, 8)),
	1071 => std_logic_vector(to_unsigned(173, 8)),
	1072 => std_logic_vector(to_unsigned(171, 8)),
	1073 => std_logic_vector(to_unsigned(168, 8)),
	1074 => std_logic_vector(to_unsigned(172, 8)),
	1075 => std_logic_vector(to_unsigned(164, 8)),
	1076 => std_logic_vector(to_unsigned(175, 8)),
	1077 => std_logic_vector(to_unsigned(168, 8)),
	1078 => std_logic_vector(to_unsigned(172, 8)),
	1079 => std_logic_vector(to_unsigned(165, 8)),
	1080 => std_logic_vector(to_unsigned(175, 8)),
	1081 => std_logic_vector(to_unsigned(170, 8)),
	1082 => std_logic_vector(to_unsigned(175, 8)),
	1083 => std_logic_vector(to_unsigned(167, 8)),
	1084 => std_logic_vector(to_unsigned(175, 8)),
	1085 => std_logic_vector(to_unsigned(165, 8)),
	1086 => std_logic_vector(to_unsigned(169, 8)),
	1087 => std_logic_vector(to_unsigned(173, 8)),
	1088 => std_logic_vector(to_unsigned(173, 8)),
	1089 => std_logic_vector(to_unsigned(162, 8)),
	1090 => std_logic_vector(to_unsigned(171, 8)),
	1091 => std_logic_vector(to_unsigned(162, 8)),
	1092 => std_logic_vector(to_unsigned(170, 8)),
	1093 => std_logic_vector(to_unsigned(163, 8)),
	1094 => std_logic_vector(to_unsigned(170, 8)),
	1095 => std_logic_vector(to_unsigned(171, 8)),
	1096 => std_logic_vector(to_unsigned(173, 8)),
	1097 => std_logic_vector(to_unsigned(169, 8)),
	1098 => std_logic_vector(to_unsigned(168, 8)),
	1099 => std_logic_vector(to_unsigned(173, 8)),
	1100 => std_logic_vector(to_unsigned(164, 8)),
	1101 => std_logic_vector(to_unsigned(171, 8)),
	1102 => std_logic_vector(to_unsigned(162, 8)),
	1103 => std_logic_vector(to_unsigned(163, 8)),
	1104 => std_logic_vector(to_unsigned(167, 8)),
	1105 => std_logic_vector(to_unsigned(173, 8)),
	1106 => std_logic_vector(to_unsigned(170, 8)),
	1107 => std_logic_vector(to_unsigned(163, 8)),
	1108 => std_logic_vector(to_unsigned(170, 8)),
	1109 => std_logic_vector(to_unsigned(165, 8)),
	1110 => std_logic_vector(to_unsigned(168, 8)),
	1111 => std_logic_vector(to_unsigned(169, 8)),
	1112 => std_logic_vector(to_unsigned(164, 8)),
	1113 => std_logic_vector(to_unsigned(163, 8)),
	1114 => std_logic_vector(to_unsigned(174, 8)),
	1115 => std_logic_vector(to_unsigned(169, 8)),
	1116 => std_logic_vector(to_unsigned(175, 8)),
	1117 => std_logic_vector(to_unsigned(176, 8)),
	1118 => std_logic_vector(to_unsigned(170, 8)),
	1119 => std_logic_vector(to_unsigned(168, 8)),
	1120 => std_logic_vector(to_unsigned(167, 8)),
	1121 => std_logic_vector(to_unsigned(163, 8)),
	1122 => std_logic_vector(to_unsigned(166, 8)),
	1123 => std_logic_vector(to_unsigned(166, 8)),
	1124 => std_logic_vector(to_unsigned(169, 8)),
	1125 => std_logic_vector(to_unsigned(172, 8)),
	1126 => std_logic_vector(to_unsigned(175, 8)),
	1127 => std_logic_vector(to_unsigned(168, 8)),
	1128 => std_logic_vector(to_unsigned(174, 8)),
	1129 => std_logic_vector(to_unsigned(162, 8)),
	1130 => std_logic_vector(to_unsigned(167, 8)),
	1131 => std_logic_vector(to_unsigned(169, 8)),
	1132 => std_logic_vector(to_unsigned(163, 8)),
	1133 => std_logic_vector(to_unsigned(173, 8)),
	1134 => std_logic_vector(to_unsigned(173, 8)),
	1135 => std_logic_vector(to_unsigned(171, 8)),
	1136 => std_logic_vector(to_unsigned(169, 8)),
	1137 => std_logic_vector(to_unsigned(173, 8)),
	1138 => std_logic_vector(to_unsigned(165, 8)),
	1139 => std_logic_vector(to_unsigned(170, 8)),
	1140 => std_logic_vector(to_unsigned(162, 8)),
	1141 => std_logic_vector(to_unsigned(170, 8)),
	1142 => std_logic_vector(to_unsigned(169, 8)),
	1143 => std_logic_vector(to_unsigned(169, 8)),
	1144 => std_logic_vector(to_unsigned(166, 8)),
	1145 => std_logic_vector(to_unsigned(174, 8)),
	1146 => std_logic_vector(to_unsigned(164, 8)),
	1147 => std_logic_vector(to_unsigned(165, 8)),
	1148 => std_logic_vector(to_unsigned(173, 8)),
	1149 => std_logic_vector(to_unsigned(173, 8)),
	1150 => std_logic_vector(to_unsigned(169, 8)),
	1151 => std_logic_vector(to_unsigned(174, 8)),
	1152 => std_logic_vector(to_unsigned(176, 8)),
	1153 => std_logic_vector(to_unsigned(172, 8)),
	1154 => std_logic_vector(to_unsigned(176, 8)),
	1155 => std_logic_vector(to_unsigned(175, 8)),
	1156 => std_logic_vector(to_unsigned(162, 8)),
	1157 => std_logic_vector(to_unsigned(166, 8)),
	1158 => std_logic_vector(to_unsigned(165, 8)),
	1159 => std_logic_vector(to_unsigned(162, 8)),
	1160 => std_logic_vector(to_unsigned(169, 8)),
	1161 => std_logic_vector(to_unsigned(175, 8)),
	1162 => std_logic_vector(to_unsigned(169, 8)),
	1163 => std_logic_vector(to_unsigned(163, 8)),
	1164 => std_logic_vector(to_unsigned(169, 8)),
	1165 => std_logic_vector(to_unsigned(162, 8)),
	1166 => std_logic_vector(to_unsigned(174, 8)),
	1167 => std_logic_vector(to_unsigned(164, 8)),
	1168 => std_logic_vector(to_unsigned(176, 8)),
	1169 => std_logic_vector(to_unsigned(163, 8)),
	1170 => std_logic_vector(to_unsigned(162, 8)),
	1171 => std_logic_vector(to_unsigned(176, 8)),
	1172 => std_logic_vector(to_unsigned(165, 8)),
	1173 => std_logic_vector(to_unsigned(168, 8)),
	1174 => std_logic_vector(to_unsigned(162, 8)),
	1175 => std_logic_vector(to_unsigned(176, 8)),
	1176 => std_logic_vector(to_unsigned(172, 8)),
	1177 => std_logic_vector(to_unsigned(169, 8)),
	1178 => std_logic_vector(to_unsigned(162, 8)),
	1179 => std_logic_vector(to_unsigned(169, 8)),
	1180 => std_logic_vector(to_unsigned(167, 8)),
	1181 => std_logic_vector(to_unsigned(172, 8)),
	1182 => std_logic_vector(to_unsigned(173, 8)),
	1183 => std_logic_vector(to_unsigned(168, 8)),
	1184 => std_logic_vector(to_unsigned(174, 8)),
	1185 => std_logic_vector(to_unsigned(164, 8)),
	1186 => std_logic_vector(to_unsigned(165, 8)),
	1187 => std_logic_vector(to_unsigned(171, 8)),
	1188 => std_logic_vector(to_unsigned(170, 8)),
	1189 => std_logic_vector(to_unsigned(175, 8)),
	1190 => std_logic_vector(to_unsigned(167, 8)),
	1191 => std_logic_vector(to_unsigned(168, 8)),
	1192 => std_logic_vector(to_unsigned(165, 8)),
	1193 => std_logic_vector(to_unsigned(165, 8)),
	1194 => std_logic_vector(to_unsigned(171, 8)),
	1195 => std_logic_vector(to_unsigned(163, 8)),
	1196 => std_logic_vector(to_unsigned(168, 8)),
	1197 => std_logic_vector(to_unsigned(168, 8)),
	1198 => std_logic_vector(to_unsigned(175, 8)),
	1199 => std_logic_vector(to_unsigned(171, 8)),
	1200 => std_logic_vector(to_unsigned(171, 8)),
	1201 => std_logic_vector(to_unsigned(166, 8)),
	1202 => std_logic_vector(to_unsigned(170, 8)),
	1203 => std_logic_vector(to_unsigned(166, 8)),
	1204 => std_logic_vector(to_unsigned(162, 8)),
	1205 => std_logic_vector(to_unsigned(172, 8)),
	1206 => std_logic_vector(to_unsigned(171, 8)),
	1207 => std_logic_vector(to_unsigned(166, 8)),
	1208 => std_logic_vector(to_unsigned(164, 8)),
	1209 => std_logic_vector(to_unsigned(163, 8)),
	1210 => std_logic_vector(to_unsigned(171, 8)),
	1211 => std_logic_vector(to_unsigned(163, 8)),
	1212 => std_logic_vector(to_unsigned(164, 8)),
	1213 => std_logic_vector(to_unsigned(163, 8)),
	1214 => std_logic_vector(to_unsigned(171, 8)),
	1215 => std_logic_vector(to_unsigned(173, 8)),
	1216 => std_logic_vector(to_unsigned(171, 8)),
	1217 => std_logic_vector(to_unsigned(176, 8)),
	1218 => std_logic_vector(to_unsigned(168, 8)),
	1219 => std_logic_vector(to_unsigned(169, 8)),
	1220 => std_logic_vector(to_unsigned(168, 8)),
	1221 => std_logic_vector(to_unsigned(176, 8)),
	1222 => std_logic_vector(to_unsigned(162, 8)),
	1223 => std_logic_vector(to_unsigned(162, 8)),
	1224 => std_logic_vector(to_unsigned(163, 8)),
	1225 => std_logic_vector(to_unsigned(171, 8)),
	1226 => std_logic_vector(to_unsigned(162, 8)),
	1227 => std_logic_vector(to_unsigned(169, 8)),
	1228 => std_logic_vector(to_unsigned(175, 8)),
	1229 => std_logic_vector(to_unsigned(162, 8)),
	1230 => std_logic_vector(to_unsigned(169, 8)),
	1231 => std_logic_vector(to_unsigned(172, 8)),
	1232 => std_logic_vector(to_unsigned(163, 8)),
	1233 => std_logic_vector(to_unsigned(175, 8)),
	1234 => std_logic_vector(to_unsigned(175, 8)),
	1235 => std_logic_vector(to_unsigned(170, 8)),
	1236 => std_logic_vector(to_unsigned(168, 8)),
	1237 => std_logic_vector(to_unsigned(176, 8)),
	1238 => std_logic_vector(to_unsigned(174, 8)),
	1239 => std_logic_vector(to_unsigned(176, 8)),
	1240 => std_logic_vector(to_unsigned(167, 8)),
	1241 => std_logic_vector(to_unsigned(167, 8)),
	1242 => std_logic_vector(to_unsigned(168, 8)),
	1243 => std_logic_vector(to_unsigned(163, 8)),
	1244 => std_logic_vector(to_unsigned(167, 8)),
	1245 => std_logic_vector(to_unsigned(170, 8)),
	1246 => std_logic_vector(to_unsigned(166, 8)),
	1247 => std_logic_vector(to_unsigned(173, 8)),
	1248 => std_logic_vector(to_unsigned(172, 8)),
	1249 => std_logic_vector(to_unsigned(176, 8)),
	1250 => std_logic_vector(to_unsigned(175, 8)),
	1251 => std_logic_vector(to_unsigned(169, 8)),
	1252 => std_logic_vector(to_unsigned(176, 8)),
	1253 => std_logic_vector(to_unsigned(164, 8)),
	1254 => std_logic_vector(to_unsigned(175, 8)),
	1255 => std_logic_vector(to_unsigned(164, 8)),
	1256 => std_logic_vector(to_unsigned(166, 8)),
	1257 => std_logic_vector(to_unsigned(165, 8)),
	1258 => std_logic_vector(to_unsigned(166, 8)),
	1259 => std_logic_vector(to_unsigned(172, 8)),
	1260 => std_logic_vector(to_unsigned(176, 8)),
	1261 => std_logic_vector(to_unsigned(170, 8)),
	1262 => std_logic_vector(to_unsigned(162, 8)),
	1263 => std_logic_vector(to_unsigned(164, 8)),
	1264 => std_logic_vector(to_unsigned(162, 8)),
	1265 => std_logic_vector(to_unsigned(165, 8)),
	1266 => std_logic_vector(to_unsigned(168, 8)),
	1267 => std_logic_vector(to_unsigned(167, 8)),
	1268 => std_logic_vector(to_unsigned(162, 8)),
	1269 => std_logic_vector(to_unsigned(171, 8)),
	1270 => std_logic_vector(to_unsigned(170, 8)),
	1271 => std_logic_vector(to_unsigned(162, 8)),
	1272 => std_logic_vector(to_unsigned(166, 8)),
	1273 => std_logic_vector(to_unsigned(175, 8)),
	1274 => std_logic_vector(to_unsigned(162, 8)),
	1275 => std_logic_vector(to_unsigned(169, 8)),
	1276 => std_logic_vector(to_unsigned(169, 8)),
	1277 => std_logic_vector(to_unsigned(174, 8)),
	1278 => std_logic_vector(to_unsigned(176, 8)),
	1279 => std_logic_vector(to_unsigned(162, 8)),
	1280 => std_logic_vector(to_unsigned(164, 8)),
	1281 => std_logic_vector(to_unsigned(174, 8)),
	1282 => std_logic_vector(to_unsigned(173, 8)),
	1283 => std_logic_vector(to_unsigned(174, 8)),
	1284 => std_logic_vector(to_unsigned(167, 8)),
	1285 => std_logic_vector(to_unsigned(163, 8)),
	1286 => std_logic_vector(to_unsigned(166, 8)),
	1287 => std_logic_vector(to_unsigned(162, 8)),
	1288 => std_logic_vector(to_unsigned(170, 8)),
	1289 => std_logic_vector(to_unsigned(166, 8)),
	1290 => std_logic_vector(to_unsigned(165, 8)),
	1291 => std_logic_vector(to_unsigned(176, 8)),
	1292 => std_logic_vector(to_unsigned(167, 8)),
	1293 => std_logic_vector(to_unsigned(173, 8)),
	1294 => std_logic_vector(to_unsigned(172, 8)),
	1295 => std_logic_vector(to_unsigned(170, 8)),
	1296 => std_logic_vector(to_unsigned(173, 8)),
	1297 => std_logic_vector(to_unsigned(165, 8)),
	1298 => std_logic_vector(to_unsigned(163, 8)),
	1299 => std_logic_vector(to_unsigned(166, 8)),
	1300 => std_logic_vector(to_unsigned(166, 8)),
	1301 => std_logic_vector(to_unsigned(168, 8)),
	1302 => std_logic_vector(to_unsigned(167, 8)),
	1303 => std_logic_vector(to_unsigned(166, 8)),
	1304 => std_logic_vector(to_unsigned(163, 8)),
	1305 => std_logic_vector(to_unsigned(175, 8)),
	1306 => std_logic_vector(to_unsigned(170, 8)),
	1307 => std_logic_vector(to_unsigned(170, 8)),
	1308 => std_logic_vector(to_unsigned(165, 8)),
	1309 => std_logic_vector(to_unsigned(162, 8)),
	1310 => std_logic_vector(to_unsigned(175, 8)),
	1311 => std_logic_vector(to_unsigned(168, 8)),
	1312 => std_logic_vector(to_unsigned(165, 8)),
	1313 => std_logic_vector(to_unsigned(172, 8)),
	1314 => std_logic_vector(to_unsigned(169, 8)),
	1315 => std_logic_vector(to_unsigned(168, 8)),
	1316 => std_logic_vector(to_unsigned(167, 8)),
	1317 => std_logic_vector(to_unsigned(171, 8)),
	1318 => std_logic_vector(to_unsigned(170, 8)),
	1319 => std_logic_vector(to_unsigned(176, 8)),
	1320 => std_logic_vector(to_unsigned(168, 8)),
	1321 => std_logic_vector(to_unsigned(169, 8)),
	1322 => std_logic_vector(to_unsigned(171, 8)),
	1323 => std_logic_vector(to_unsigned(174, 8)),
	1324 => std_logic_vector(to_unsigned(167, 8)),
	1325 => std_logic_vector(to_unsigned(175, 8)),
	1326 => std_logic_vector(to_unsigned(173, 8)),
	1327 => std_logic_vector(to_unsigned(173, 8)),
	1328 => std_logic_vector(to_unsigned(167, 8)),
	1329 => std_logic_vector(to_unsigned(164, 8)),
	1330 => std_logic_vector(to_unsigned(174, 8)),
	1331 => std_logic_vector(to_unsigned(166, 8)),
	1332 => std_logic_vector(to_unsigned(171, 8)),
	1333 => std_logic_vector(to_unsigned(174, 8)),
	1334 => std_logic_vector(to_unsigned(173, 8)),
	1335 => std_logic_vector(to_unsigned(165, 8)),
	1336 => std_logic_vector(to_unsigned(164, 8)),
	1337 => std_logic_vector(to_unsigned(163, 8)),
	1338 => std_logic_vector(to_unsigned(166, 8)),
	1339 => std_logic_vector(to_unsigned(174, 8)),
	1340 => std_logic_vector(to_unsigned(176, 8)),
	1341 => std_logic_vector(to_unsigned(173, 8)),
	1342 => std_logic_vector(to_unsigned(168, 8)),
	1343 => std_logic_vector(to_unsigned(176, 8)),
	1344 => std_logic_vector(to_unsigned(168, 8)),
	1345 => std_logic_vector(to_unsigned(172, 8)),
	1346 => std_logic_vector(to_unsigned(168, 8)),
	1347 => std_logic_vector(to_unsigned(171, 8)),
	1348 => std_logic_vector(to_unsigned(172, 8)),
	1349 => std_logic_vector(to_unsigned(174, 8)),
	1350 => std_logic_vector(to_unsigned(166, 8)),
	1351 => std_logic_vector(to_unsigned(173, 8)),
	1352 => std_logic_vector(to_unsigned(170, 8)),
	1353 => std_logic_vector(to_unsigned(167, 8)),
	1354 => std_logic_vector(to_unsigned(171, 8)),
	1355 => std_logic_vector(to_unsigned(166, 8)),
	1356 => std_logic_vector(to_unsigned(175, 8)),
	1357 => std_logic_vector(to_unsigned(162, 8)),
	1358 => std_logic_vector(to_unsigned(168, 8)),
	1359 => std_logic_vector(to_unsigned(167, 8)),
	1360 => std_logic_vector(to_unsigned(172, 8)),
	1361 => std_logic_vector(to_unsigned(168, 8)),
	1362 => std_logic_vector(to_unsigned(171, 8)),
	1363 => std_logic_vector(to_unsigned(176, 8)),
	1364 => std_logic_vector(to_unsigned(164, 8)),
	1365 => std_logic_vector(to_unsigned(167, 8)),
	1366 => std_logic_vector(to_unsigned(175, 8)),
	1367 => std_logic_vector(to_unsigned(170, 8)),
	1368 => std_logic_vector(to_unsigned(173, 8)),
	1369 => std_logic_vector(to_unsigned(166, 8)),
	1370 => std_logic_vector(to_unsigned(172, 8)),
	1371 => std_logic_vector(to_unsigned(173, 8)),
	1372 => std_logic_vector(to_unsigned(167, 8)),
	1373 => std_logic_vector(to_unsigned(163, 8)),
	1374 => std_logic_vector(to_unsigned(175, 8)),
	1375 => std_logic_vector(to_unsigned(166, 8)),
	1376 => std_logic_vector(to_unsigned(168, 8)),
	1377 => std_logic_vector(to_unsigned(173, 8)),
	1378 => std_logic_vector(to_unsigned(174, 8)),
	1379 => std_logic_vector(to_unsigned(162, 8)),
	1380 => std_logic_vector(to_unsigned(173, 8)),
	1381 => std_logic_vector(to_unsigned(162, 8)),
	1382 => std_logic_vector(to_unsigned(171, 8)),
	1383 => std_logic_vector(to_unsigned(172, 8)),
	1384 => std_logic_vector(to_unsigned(169, 8)),
	1385 => std_logic_vector(to_unsigned(170, 8)),
	1386 => std_logic_vector(to_unsigned(176, 8)),
	1387 => std_logic_vector(to_unsigned(172, 8)),
	1388 => std_logic_vector(to_unsigned(176, 8)),
	1389 => std_logic_vector(to_unsigned(164, 8)),
	1390 => std_logic_vector(to_unsigned(167, 8)),
	1391 => std_logic_vector(to_unsigned(176, 8)),
	1392 => std_logic_vector(to_unsigned(164, 8)),
	1393 => std_logic_vector(to_unsigned(176, 8)),
	1394 => std_logic_vector(to_unsigned(170, 8)),
	1395 => std_logic_vector(to_unsigned(166, 8)),
	1396 => std_logic_vector(to_unsigned(171, 8)),
	1397 => std_logic_vector(to_unsigned(175, 8)),
	1398 => std_logic_vector(to_unsigned(168, 8)),
	1399 => std_logic_vector(to_unsigned(166, 8)),
	1400 => std_logic_vector(to_unsigned(173, 8)),
	1401 => std_logic_vector(to_unsigned(163, 8)),
	1402 => std_logic_vector(to_unsigned(164, 8)),
	1403 => std_logic_vector(to_unsigned(170, 8)),
	1404 => std_logic_vector(to_unsigned(165, 8)),
	1405 => std_logic_vector(to_unsigned(165, 8)),
	1406 => std_logic_vector(to_unsigned(174, 8)),
	1407 => std_logic_vector(to_unsigned(176, 8)),
	1408 => std_logic_vector(to_unsigned(172, 8)),
	1409 => std_logic_vector(to_unsigned(164, 8)),
	1410 => std_logic_vector(to_unsigned(166, 8)),
	1411 => std_logic_vector(to_unsigned(167, 8)),
	1412 => std_logic_vector(to_unsigned(174, 8)),
	1413 => std_logic_vector(to_unsigned(165, 8)),
	1414 => std_logic_vector(to_unsigned(163, 8)),
	1415 => std_logic_vector(to_unsigned(176, 8)),
	1416 => std_logic_vector(to_unsigned(176, 8)),
	1417 => std_logic_vector(to_unsigned(162, 8)),
	1418 => std_logic_vector(to_unsigned(170, 8)),
	1419 => std_logic_vector(to_unsigned(169, 8)),
	1420 => std_logic_vector(to_unsigned(168, 8)),
	1421 => std_logic_vector(to_unsigned(164, 8)),
	1422 => std_logic_vector(to_unsigned(168, 8)),
	1423 => std_logic_vector(to_unsigned(170, 8)),
	1424 => std_logic_vector(to_unsigned(172, 8)),
	1425 => std_logic_vector(to_unsigned(174, 8)),
	1426 => std_logic_vector(to_unsigned(166, 8)),
	1427 => std_logic_vector(to_unsigned(176, 8)),
	1428 => std_logic_vector(to_unsigned(167, 8)),
	1429 => std_logic_vector(to_unsigned(162, 8)),
	1430 => std_logic_vector(to_unsigned(169, 8)),
	1431 => std_logic_vector(to_unsigned(166, 8)),
	1432 => std_logic_vector(to_unsigned(175, 8)),
	1433 => std_logic_vector(to_unsigned(176, 8)),
	1434 => std_logic_vector(to_unsigned(176, 8)),
	1435 => std_logic_vector(to_unsigned(167, 8)),
	1436 => std_logic_vector(to_unsigned(176, 8)),
	1437 => std_logic_vector(to_unsigned(176, 8)),
	1438 => std_logic_vector(to_unsigned(176, 8)),
	1439 => std_logic_vector(to_unsigned(162, 8)),
	1440 => std_logic_vector(to_unsigned(162, 8)),
	1441 => std_logic_vector(to_unsigned(176, 8)),
	1442 => std_logic_vector(to_unsigned(169, 8)),
	1443 => std_logic_vector(to_unsigned(163, 8)),
	1444 => std_logic_vector(to_unsigned(171, 8)),
	1445 => std_logic_vector(to_unsigned(167, 8)),
	1446 => std_logic_vector(to_unsigned(171, 8)),
	1447 => std_logic_vector(to_unsigned(162, 8)),
	1448 => std_logic_vector(to_unsigned(173, 8)),
	1449 => std_logic_vector(to_unsigned(165, 8)),
	1450 => std_logic_vector(to_unsigned(166, 8)),
	1451 => std_logic_vector(to_unsigned(162, 8)),
	1452 => std_logic_vector(to_unsigned(176, 8)),
	1453 => std_logic_vector(to_unsigned(164, 8)),
	1454 => std_logic_vector(to_unsigned(163, 8)),
	1455 => std_logic_vector(to_unsigned(162, 8)),
	1456 => std_logic_vector(to_unsigned(173, 8)),
	1457 => std_logic_vector(to_unsigned(176, 8)),
	1458 => std_logic_vector(to_unsigned(175, 8)),
	1459 => std_logic_vector(to_unsigned(176, 8)),
	1460 => std_logic_vector(to_unsigned(168, 8)),
	1461 => std_logic_vector(to_unsigned(167, 8)),
	1462 => std_logic_vector(to_unsigned(170, 8)),
	1463 => std_logic_vector(to_unsigned(174, 8)),
	1464 => std_logic_vector(to_unsigned(162, 8)),
	1465 => std_logic_vector(to_unsigned(166, 8)),
	1466 => std_logic_vector(to_unsigned(173, 8)),
	1467 => std_logic_vector(to_unsigned(168, 8)),
	1468 => std_logic_vector(to_unsigned(168, 8)),
	1469 => std_logic_vector(to_unsigned(169, 8)),
	1470 => std_logic_vector(to_unsigned(173, 8)),
	1471 => std_logic_vector(to_unsigned(174, 8)),
	1472 => std_logic_vector(to_unsigned(162, 8)),
	1473 => std_logic_vector(to_unsigned(175, 8)),
	1474 => std_logic_vector(to_unsigned(170, 8)),
	1475 => std_logic_vector(to_unsigned(172, 8)),
	1476 => std_logic_vector(to_unsigned(169, 8)),
	1477 => std_logic_vector(to_unsigned(175, 8)),
	1478 => std_logic_vector(to_unsigned(170, 8)),
	1479 => std_logic_vector(to_unsigned(167, 8)),
	1480 => std_logic_vector(to_unsigned(163, 8)),
	1481 => std_logic_vector(to_unsigned(167, 8)),
	1482 => std_logic_vector(to_unsigned(165, 8)),
	1483 => std_logic_vector(to_unsigned(173, 8)),
	1484 => std_logic_vector(to_unsigned(169, 8)),
	1485 => std_logic_vector(to_unsigned(175, 8)),
	1486 => std_logic_vector(to_unsigned(171, 8)),
	1487 => std_logic_vector(to_unsigned(162, 8)),
	1488 => std_logic_vector(to_unsigned(174, 8)),
	1489 => std_logic_vector(to_unsigned(167, 8)),
	1490 => std_logic_vector(to_unsigned(163, 8)),
	1491 => std_logic_vector(to_unsigned(169, 8)),
	1492 => std_logic_vector(to_unsigned(170, 8)),
	1493 => std_logic_vector(to_unsigned(176, 8)),
	1494 => std_logic_vector(to_unsigned(165, 8)),
	1495 => std_logic_vector(to_unsigned(169, 8)),
	1496 => std_logic_vector(to_unsigned(170, 8)),
	1497 => std_logic_vector(to_unsigned(173, 8)),
	1498 => std_logic_vector(to_unsigned(167, 8)),
	1499 => std_logic_vector(to_unsigned(162, 8)),
	1500 => std_logic_vector(to_unsigned(168, 8)),
	1501 => std_logic_vector(to_unsigned(171, 8)),
	1502 => std_logic_vector(to_unsigned(163, 8)),
	1503 => std_logic_vector(to_unsigned(171, 8)),
	1504 => std_logic_vector(to_unsigned(171, 8)),
	1505 => std_logic_vector(to_unsigned(166, 8)),
	1506 => std_logic_vector(to_unsigned(168, 8)),
	1507 => std_logic_vector(to_unsigned(166, 8)),
	1508 => std_logic_vector(to_unsigned(172, 8)),
	1509 => std_logic_vector(to_unsigned(165, 8)),
	1510 => std_logic_vector(to_unsigned(173, 8)),
	1511 => std_logic_vector(to_unsigned(165, 8)),
	1512 => std_logic_vector(to_unsigned(173, 8)),
	1513 => std_logic_vector(to_unsigned(168, 8)),
	1514 => std_logic_vector(to_unsigned(176, 8)),
	1515 => std_logic_vector(to_unsigned(176, 8)),
	1516 => std_logic_vector(to_unsigned(171, 8)),
	1517 => std_logic_vector(to_unsigned(165, 8)),
	1518 => std_logic_vector(to_unsigned(170, 8)),
	1519 => std_logic_vector(to_unsigned(168, 8)),
	1520 => std_logic_vector(to_unsigned(172, 8)),
	1521 => std_logic_vector(to_unsigned(175, 8)),
	1522 => std_logic_vector(to_unsigned(173, 8)),
	1523 => std_logic_vector(to_unsigned(165, 8)),
	1524 => std_logic_vector(to_unsigned(171, 8)),
	1525 => std_logic_vector(to_unsigned(172, 8)),
	1526 => std_logic_vector(to_unsigned(165, 8)),
	1527 => std_logic_vector(to_unsigned(163, 8)),
	1528 => std_logic_vector(to_unsigned(175, 8)),
	1529 => std_logic_vector(to_unsigned(175, 8)),
	1530 => std_logic_vector(to_unsigned(165, 8)),
	1531 => std_logic_vector(to_unsigned(172, 8)),
	1532 => std_logic_vector(to_unsigned(162, 8)),
	1533 => std_logic_vector(to_unsigned(162, 8)),
	1534 => std_logic_vector(to_unsigned(173, 8)),
	1535 => std_logic_vector(to_unsigned(167, 8)),
	1536 => std_logic_vector(to_unsigned(176, 8)),
	1537 => std_logic_vector(to_unsigned(175, 8)),
	1538 => std_logic_vector(to_unsigned(175, 8)),
	1539 => std_logic_vector(to_unsigned(168, 8)),
	1540 => std_logic_vector(to_unsigned(170, 8)),
	1541 => std_logic_vector(to_unsigned(169, 8)),
	1542 => std_logic_vector(to_unsigned(167, 8)),
	1543 => std_logic_vector(to_unsigned(174, 8)),
	1544 => std_logic_vector(to_unsigned(168, 8)),
	1545 => std_logic_vector(to_unsigned(165, 8)),
	1546 => std_logic_vector(to_unsigned(164, 8)),
	1547 => std_logic_vector(to_unsigned(174, 8)),
	1548 => std_logic_vector(to_unsigned(167, 8)),
	1549 => std_logic_vector(to_unsigned(166, 8)),
	1550 => std_logic_vector(to_unsigned(163, 8)),
	1551 => std_logic_vector(to_unsigned(175, 8)),
	1552 => std_logic_vector(to_unsigned(172, 8)),
	1553 => std_logic_vector(to_unsigned(175, 8)),
	1554 => std_logic_vector(to_unsigned(166, 8)),
	1555 => std_logic_vector(to_unsigned(170, 8)),
	1556 => std_logic_vector(to_unsigned(163, 8)),
	1557 => std_logic_vector(to_unsigned(172, 8)),
	1558 => std_logic_vector(to_unsigned(176, 8)),
	1559 => std_logic_vector(to_unsigned(164, 8)),
	1560 => std_logic_vector(to_unsigned(169, 8)),
	1561 => std_logic_vector(to_unsigned(162, 8)),
	1562 => std_logic_vector(to_unsigned(173, 8)),
	1563 => std_logic_vector(to_unsigned(176, 8)),
	1564 => std_logic_vector(to_unsigned(171, 8)),
	1565 => std_logic_vector(to_unsigned(164, 8)),
	1566 => std_logic_vector(to_unsigned(163, 8)),
	1567 => std_logic_vector(to_unsigned(170, 8)),
	1568 => std_logic_vector(to_unsigned(165, 8)),
	1569 => std_logic_vector(to_unsigned(164, 8)),
	1570 => std_logic_vector(to_unsigned(164, 8)),
	1571 => std_logic_vector(to_unsigned(163, 8)),
	1572 => std_logic_vector(to_unsigned(164, 8)),
	1573 => std_logic_vector(to_unsigned(172, 8)),
	1574 => std_logic_vector(to_unsigned(171, 8)),
	1575 => std_logic_vector(to_unsigned(176, 8)),
	1576 => std_logic_vector(to_unsigned(167, 8)),
	1577 => std_logic_vector(to_unsigned(175, 8)),
	1578 => std_logic_vector(to_unsigned(164, 8)),
	1579 => std_logic_vector(to_unsigned(172, 8)),
	1580 => std_logic_vector(to_unsigned(170, 8)),
	1581 => std_logic_vector(to_unsigned(163, 8)),
	1582 => std_logic_vector(to_unsigned(172, 8)),
	1583 => std_logic_vector(to_unsigned(170, 8)),
	1584 => std_logic_vector(to_unsigned(176, 8)),
	1585 => std_logic_vector(to_unsigned(163, 8)),
	1586 => std_logic_vector(to_unsigned(171, 8)),
	1587 => std_logic_vector(to_unsigned(165, 8)),
	1588 => std_logic_vector(to_unsigned(165, 8)),
	1589 => std_logic_vector(to_unsigned(170, 8)),
	1590 => std_logic_vector(to_unsigned(168, 8)),
	1591 => std_logic_vector(to_unsigned(170, 8)),
	1592 => std_logic_vector(to_unsigned(167, 8)),
	1593 => std_logic_vector(to_unsigned(162, 8)),
	1594 => std_logic_vector(to_unsigned(168, 8)),
	1595 => std_logic_vector(to_unsigned(176, 8)),
	1596 => std_logic_vector(to_unsigned(172, 8)),
	1597 => std_logic_vector(to_unsigned(168, 8)),
	1598 => std_logic_vector(to_unsigned(170, 8)),
	1599 => std_logic_vector(to_unsigned(172, 8)),
	1600 => std_logic_vector(to_unsigned(168, 8)),
	1601 => std_logic_vector(to_unsigned(163, 8)),
	1602 => std_logic_vector(to_unsigned(169, 8)),
	1603 => std_logic_vector(to_unsigned(163, 8)),
	1604 => std_logic_vector(to_unsigned(176, 8)),
	1605 => std_logic_vector(to_unsigned(175, 8)),
	1606 => std_logic_vector(to_unsigned(171, 8)),
	1607 => std_logic_vector(to_unsigned(167, 8)),
	1608 => std_logic_vector(to_unsigned(162, 8)),
	1609 => std_logic_vector(to_unsigned(174, 8)),
	1610 => std_logic_vector(to_unsigned(167, 8)),
	1611 => std_logic_vector(to_unsigned(166, 8)),
	1612 => std_logic_vector(to_unsigned(174, 8)),
	1613 => std_logic_vector(to_unsigned(176, 8)),
	1614 => std_logic_vector(to_unsigned(173, 8)),
	1615 => std_logic_vector(to_unsigned(167, 8)),
	1616 => std_logic_vector(to_unsigned(171, 8)),
	1617 => std_logic_vector(to_unsigned(171, 8)),
	1618 => std_logic_vector(to_unsigned(171, 8)),
	1619 => std_logic_vector(to_unsigned(170, 8)),
	1620 => std_logic_vector(to_unsigned(167, 8)),
	1621 => std_logic_vector(to_unsigned(173, 8)),
	1622 => std_logic_vector(to_unsigned(162, 8)),
	1623 => std_logic_vector(to_unsigned(167, 8)),
	1624 => std_logic_vector(to_unsigned(167, 8)),
	1625 => std_logic_vector(to_unsigned(171, 8)),
	1626 => std_logic_vector(to_unsigned(166, 8)),
	1627 => std_logic_vector(to_unsigned(172, 8)),
	1628 => std_logic_vector(to_unsigned(163, 8)),
	1629 => std_logic_vector(to_unsigned(172, 8)),
	1630 => std_logic_vector(to_unsigned(172, 8)),
	1631 => std_logic_vector(to_unsigned(174, 8)),
	1632 => std_logic_vector(to_unsigned(171, 8)),
	1633 => std_logic_vector(to_unsigned(172, 8)),
	1634 => std_logic_vector(to_unsigned(171, 8)),
	1635 => std_logic_vector(to_unsigned(170, 8)),
	1636 => std_logic_vector(to_unsigned(164, 8)),
	1637 => std_logic_vector(to_unsigned(162, 8)),
	1638 => std_logic_vector(to_unsigned(170, 8)),
	1639 => std_logic_vector(to_unsigned(171, 8)),
	1640 => std_logic_vector(to_unsigned(162, 8)),
	1641 => std_logic_vector(to_unsigned(174, 8)),
	1642 => std_logic_vector(to_unsigned(171, 8)),
	1643 => std_logic_vector(to_unsigned(171, 8)),
	1644 => std_logic_vector(to_unsigned(176, 8)),
	1645 => std_logic_vector(to_unsigned(173, 8)),
	1646 => std_logic_vector(to_unsigned(175, 8)),
	1647 => std_logic_vector(to_unsigned(171, 8)),
	1648 => std_logic_vector(to_unsigned(166, 8)),
	1649 => std_logic_vector(to_unsigned(168, 8)),
	1650 => std_logic_vector(to_unsigned(173, 8)),
	1651 => std_logic_vector(to_unsigned(163, 8)),
	1652 => std_logic_vector(to_unsigned(175, 8)),
	1653 => std_logic_vector(to_unsigned(166, 8)),
	1654 => std_logic_vector(to_unsigned(165, 8)),
	1655 => std_logic_vector(to_unsigned(169, 8)),
	1656 => std_logic_vector(to_unsigned(163, 8)),
	1657 => std_logic_vector(to_unsigned(165, 8)),
	1658 => std_logic_vector(to_unsigned(163, 8)),
	1659 => std_logic_vector(to_unsigned(175, 8)),
	1660 => std_logic_vector(to_unsigned(167, 8)),
	1661 => std_logic_vector(to_unsigned(174, 8)),
	1662 => std_logic_vector(to_unsigned(167, 8)),
	1663 => std_logic_vector(to_unsigned(164, 8)),
	1664 => std_logic_vector(to_unsigned(173, 8)),
	1665 => std_logic_vector(to_unsigned(171, 8)),
	1666 => std_logic_vector(to_unsigned(170, 8)),
	1667 => std_logic_vector(to_unsigned(169, 8)),
	1668 => std_logic_vector(to_unsigned(164, 8)),
	1669 => std_logic_vector(to_unsigned(169, 8)),
	1670 => std_logic_vector(to_unsigned(171, 8)),
	1671 => std_logic_vector(to_unsigned(173, 8)),
	1672 => std_logic_vector(to_unsigned(170, 8)),
	1673 => std_logic_vector(to_unsigned(176, 8)),
	1674 => std_logic_vector(to_unsigned(169, 8)),
	1675 => std_logic_vector(to_unsigned(171, 8)),
	1676 => std_logic_vector(to_unsigned(163, 8)),
	1677 => std_logic_vector(to_unsigned(173, 8)),
	1678 => std_logic_vector(to_unsigned(173, 8)),
	1679 => std_logic_vector(to_unsigned(171, 8)),
	1680 => std_logic_vector(to_unsigned(169, 8)),
	1681 => std_logic_vector(to_unsigned(173, 8)),
	1682 => std_logic_vector(to_unsigned(169, 8)),
	1683 => std_logic_vector(to_unsigned(175, 8)),
	1684 => std_logic_vector(to_unsigned(164, 8)),
	1685 => std_logic_vector(to_unsigned(175, 8)),
	1686 => std_logic_vector(to_unsigned(166, 8)),
	1687 => std_logic_vector(to_unsigned(164, 8)),
	1688 => std_logic_vector(to_unsigned(163, 8)),
	1689 => std_logic_vector(to_unsigned(162, 8)),
	1690 => std_logic_vector(to_unsigned(170, 8)),
	1691 => std_logic_vector(to_unsigned(175, 8)),
	1692 => std_logic_vector(to_unsigned(168, 8)),
	1693 => std_logic_vector(to_unsigned(176, 8)),
	1694 => std_logic_vector(to_unsigned(170, 8)),
	1695 => std_logic_vector(to_unsigned(172, 8)),
	1696 => std_logic_vector(to_unsigned(165, 8)),
	1697 => std_logic_vector(to_unsigned(167, 8)),
	1698 => std_logic_vector(to_unsigned(171, 8)),
	1699 => std_logic_vector(to_unsigned(166, 8)),
	1700 => std_logic_vector(to_unsigned(173, 8)),
	1701 => std_logic_vector(to_unsigned(163, 8)),
	1702 => std_logic_vector(to_unsigned(166, 8)),
	1703 => std_logic_vector(to_unsigned(172, 8)),
	1704 => std_logic_vector(to_unsigned(168, 8)),
	1705 => std_logic_vector(to_unsigned(162, 8)),
	1706 => std_logic_vector(to_unsigned(174, 8)),
	1707 => std_logic_vector(to_unsigned(167, 8)),
	1708 => std_logic_vector(to_unsigned(164, 8)),
	1709 => std_logic_vector(to_unsigned(175, 8)),
	1710 => std_logic_vector(to_unsigned(169, 8)),
	1711 => std_logic_vector(to_unsigned(164, 8)),
	1712 => std_logic_vector(to_unsigned(175, 8)),
	1713 => std_logic_vector(to_unsigned(171, 8)),
	1714 => std_logic_vector(to_unsigned(165, 8)),
	1715 => std_logic_vector(to_unsigned(172, 8)),
	1716 => std_logic_vector(to_unsigned(166, 8)),
	1717 => std_logic_vector(to_unsigned(165, 8)),
	1718 => std_logic_vector(to_unsigned(174, 8)),
	1719 => std_logic_vector(to_unsigned(165, 8)),
	1720 => std_logic_vector(to_unsigned(167, 8)),
	1721 => std_logic_vector(to_unsigned(162, 8)),
	1722 => std_logic_vector(to_unsigned(175, 8)),
	1723 => std_logic_vector(to_unsigned(174, 8)),
	1724 => std_logic_vector(to_unsigned(165, 8)),
	1725 => std_logic_vector(to_unsigned(173, 8)),
	1726 => std_logic_vector(to_unsigned(165, 8)),
	1727 => std_logic_vector(to_unsigned(173, 8)),
	1728 => std_logic_vector(to_unsigned(169, 8)),
	1729 => std_logic_vector(to_unsigned(165, 8)),
	1730 => std_logic_vector(to_unsigned(171, 8)),
	1731 => std_logic_vector(to_unsigned(164, 8)),
	1732 => std_logic_vector(to_unsigned(166, 8)),
	1733 => std_logic_vector(to_unsigned(175, 8)),
	1734 => std_logic_vector(to_unsigned(168, 8)),
	1735 => std_logic_vector(to_unsigned(167, 8)),
	1736 => std_logic_vector(to_unsigned(174, 8)),
	1737 => std_logic_vector(to_unsigned(167, 8)),
	1738 => std_logic_vector(to_unsigned(163, 8)),
	1739 => std_logic_vector(to_unsigned(162, 8)),
	1740 => std_logic_vector(to_unsigned(169, 8)),
	1741 => std_logic_vector(to_unsigned(170, 8)),
	1742 => std_logic_vector(to_unsigned(164, 8)),
	1743 => std_logic_vector(to_unsigned(163, 8)),
	1744 => std_logic_vector(to_unsigned(176, 8)),
	1745 => std_logic_vector(to_unsigned(165, 8)),
	1746 => std_logic_vector(to_unsigned(175, 8)),
	1747 => std_logic_vector(to_unsigned(175, 8)),
	1748 => std_logic_vector(to_unsigned(165, 8)),
	1749 => std_logic_vector(to_unsigned(164, 8)),
	1750 => std_logic_vector(to_unsigned(171, 8)),
	1751 => std_logic_vector(to_unsigned(176, 8)),
	1752 => std_logic_vector(to_unsigned(174, 8)),
	1753 => std_logic_vector(to_unsigned(162, 8)),
	1754 => std_logic_vector(to_unsigned(170, 8)),
	1755 => std_logic_vector(to_unsigned(173, 8)),
	1756 => std_logic_vector(to_unsigned(167, 8)),
	1757 => std_logic_vector(to_unsigned(162, 8)),
	1758 => std_logic_vector(to_unsigned(176, 8)),
	1759 => std_logic_vector(to_unsigned(167, 8)),
	1760 => std_logic_vector(to_unsigned(167, 8)),
	1761 => std_logic_vector(to_unsigned(169, 8)),
	1762 => std_logic_vector(to_unsigned(165, 8)),
	1763 => std_logic_vector(to_unsigned(176, 8)),
	1764 => std_logic_vector(to_unsigned(169, 8)),
	1765 => std_logic_vector(to_unsigned(166, 8)),
	1766 => std_logic_vector(to_unsigned(167, 8)),
	1767 => std_logic_vector(to_unsigned(166, 8)),
	1768 => std_logic_vector(to_unsigned(175, 8)),
	1769 => std_logic_vector(to_unsigned(174, 8)),
	1770 => std_logic_vector(to_unsigned(175, 8)),
	1771 => std_logic_vector(to_unsigned(166, 8)),
	1772 => std_logic_vector(to_unsigned(171, 8)),
	1773 => std_logic_vector(to_unsigned(165, 8)),
	1774 => std_logic_vector(to_unsigned(169, 8)),
	1775 => std_logic_vector(to_unsigned(173, 8)),
	1776 => std_logic_vector(to_unsigned(166, 8)),
	1777 => std_logic_vector(to_unsigned(167, 8)),
	1778 => std_logic_vector(to_unsigned(165, 8)),
	1779 => std_logic_vector(to_unsigned(174, 8)),
	1780 => std_logic_vector(to_unsigned(171, 8)),
	1781 => std_logic_vector(to_unsigned(164, 8)),
	1782 => std_logic_vector(to_unsigned(164, 8)),
	1783 => std_logic_vector(to_unsigned(171, 8)),
	1784 => std_logic_vector(to_unsigned(170, 8)),
	1785 => std_logic_vector(to_unsigned(171, 8)),
	1786 => std_logic_vector(to_unsigned(172, 8)),
	1787 => std_logic_vector(to_unsigned(171, 8)),
	1788 => std_logic_vector(to_unsigned(162, 8)),
	1789 => std_logic_vector(to_unsigned(169, 8)),
	1790 => std_logic_vector(to_unsigned(176, 8)),
	1791 => std_logic_vector(to_unsigned(165, 8)),
	1792 => std_logic_vector(to_unsigned(171, 8)),
	1793 => std_logic_vector(to_unsigned(173, 8)),
	1794 => std_logic_vector(to_unsigned(175, 8)),
	1795 => std_logic_vector(to_unsigned(175, 8)),
	1796 => std_logic_vector(to_unsigned(175, 8)),
	1797 => std_logic_vector(to_unsigned(174, 8)),
	1798 => std_logic_vector(to_unsigned(164, 8)),
	1799 => std_logic_vector(to_unsigned(175, 8)),
	1800 => std_logic_vector(to_unsigned(171, 8)),
	1801 => std_logic_vector(to_unsigned(171, 8)),
	1802 => std_logic_vector(to_unsigned(174, 8)),
	1803 => std_logic_vector(to_unsigned(172, 8)),
	1804 => std_logic_vector(to_unsigned(162, 8)),
	1805 => std_logic_vector(to_unsigned(172, 8)),
	1806 => std_logic_vector(to_unsigned(167, 8)),
	1807 => std_logic_vector(to_unsigned(174, 8)),
	1808 => std_logic_vector(to_unsigned(172, 8)),
	1809 => std_logic_vector(to_unsigned(166, 8)),
	1810 => std_logic_vector(to_unsigned(170, 8)),
	1811 => std_logic_vector(to_unsigned(170, 8)),
	1812 => std_logic_vector(to_unsigned(175, 8)),
	1813 => std_logic_vector(to_unsigned(165, 8)),
	1814 => std_logic_vector(to_unsigned(169, 8)),
	1815 => std_logic_vector(to_unsigned(166, 8)),
	1816 => std_logic_vector(to_unsigned(164, 8)),
	1817 => std_logic_vector(to_unsigned(169, 8)),
	1818 => std_logic_vector(to_unsigned(168, 8)),
	1819 => std_logic_vector(to_unsigned(171, 8)),
	1820 => std_logic_vector(to_unsigned(169, 8)),
	1821 => std_logic_vector(to_unsigned(172, 8)),
	1822 => std_logic_vector(to_unsigned(176, 8)),
	1823 => std_logic_vector(to_unsigned(165, 8)),
	1824 => std_logic_vector(to_unsigned(163, 8)),
	1825 => std_logic_vector(to_unsigned(165, 8)),
	1826 => std_logic_vector(to_unsigned(164, 8)),
	1827 => std_logic_vector(to_unsigned(176, 8)),
	1828 => std_logic_vector(to_unsigned(171, 8)),
	1829 => std_logic_vector(to_unsigned(171, 8)),
	1830 => std_logic_vector(to_unsigned(168, 8)),
	1831 => std_logic_vector(to_unsigned(173, 8)),
	1832 => std_logic_vector(to_unsigned(167, 8)),
	1833 => std_logic_vector(to_unsigned(166, 8)),
	1834 => std_logic_vector(to_unsigned(174, 8)),
	1835 => std_logic_vector(to_unsigned(165, 8)),
	1836 => std_logic_vector(to_unsigned(170, 8)),
	1837 => std_logic_vector(to_unsigned(162, 8)),
	1838 => std_logic_vector(to_unsigned(169, 8)),
	1839 => std_logic_vector(to_unsigned(167, 8)),
	1840 => std_logic_vector(to_unsigned(166, 8)),
	1841 => std_logic_vector(to_unsigned(176, 8)),
	1842 => std_logic_vector(to_unsigned(168, 8)),
	1843 => std_logic_vector(to_unsigned(169, 8)),
	1844 => std_logic_vector(to_unsigned(165, 8)),
	1845 => std_logic_vector(to_unsigned(169, 8)),
	1846 => std_logic_vector(to_unsigned(175, 8)),
	1847 => std_logic_vector(to_unsigned(166, 8)),
	1848 => std_logic_vector(to_unsigned(169, 8)),
	1849 => std_logic_vector(to_unsigned(171, 8)),
	1850 => std_logic_vector(to_unsigned(174, 8)),
	1851 => std_logic_vector(to_unsigned(167, 8)),
	1852 => std_logic_vector(to_unsigned(162, 8)),
	1853 => std_logic_vector(to_unsigned(175, 8)),
	1854 => std_logic_vector(to_unsigned(174, 8)),
	1855 => std_logic_vector(to_unsigned(174, 8)),
	1856 => std_logic_vector(to_unsigned(168, 8)),
	1857 => std_logic_vector(to_unsigned(173, 8)),
	1858 => std_logic_vector(to_unsigned(163, 8)),
	1859 => std_logic_vector(to_unsigned(176, 8)),
	1860 => std_logic_vector(to_unsigned(170, 8)),
	1861 => std_logic_vector(to_unsigned(172, 8)),
	1862 => std_logic_vector(to_unsigned(168, 8)),
	1863 => std_logic_vector(to_unsigned(162, 8)),
	1864 => std_logic_vector(to_unsigned(173, 8)),
	1865 => std_logic_vector(to_unsigned(175, 8)),
	1866 => std_logic_vector(to_unsigned(172, 8)),
	1867 => std_logic_vector(to_unsigned(175, 8)),
	1868 => std_logic_vector(to_unsigned(174, 8)),
	1869 => std_logic_vector(to_unsigned(174, 8)),
	1870 => std_logic_vector(to_unsigned(169, 8)),
	1871 => std_logic_vector(to_unsigned(176, 8)),
	1872 => std_logic_vector(to_unsigned(164, 8)),
	1873 => std_logic_vector(to_unsigned(170, 8)),
	1874 => std_logic_vector(to_unsigned(175, 8)),
	1875 => std_logic_vector(to_unsigned(170, 8)),
	1876 => std_logic_vector(to_unsigned(162, 8)),
	1877 => std_logic_vector(to_unsigned(172, 8)),
	1878 => std_logic_vector(to_unsigned(166, 8)),
	1879 => std_logic_vector(to_unsigned(173, 8)),
	1880 => std_logic_vector(to_unsigned(174, 8)),
	1881 => std_logic_vector(to_unsigned(172, 8)),
	1882 => std_logic_vector(to_unsigned(173, 8)),
	1883 => std_logic_vector(to_unsigned(165, 8)),
	1884 => std_logic_vector(to_unsigned(162, 8)),
	1885 => std_logic_vector(to_unsigned(175, 8)),
	1886 => std_logic_vector(to_unsigned(176, 8)),
	1887 => std_logic_vector(to_unsigned(170, 8)),
	1888 => std_logic_vector(to_unsigned(165, 8)),
	1889 => std_logic_vector(to_unsigned(171, 8)),
	1890 => std_logic_vector(to_unsigned(169, 8)),
	1891 => std_logic_vector(to_unsigned(166, 8)),
	1892 => std_logic_vector(to_unsigned(163, 8)),
	1893 => std_logic_vector(to_unsigned(170, 8)),
	1894 => std_logic_vector(to_unsigned(170, 8)),
	1895 => std_logic_vector(to_unsigned(168, 8)),
	1896 => std_logic_vector(to_unsigned(171, 8)),
	1897 => std_logic_vector(to_unsigned(176, 8)),
	1898 => std_logic_vector(to_unsigned(167, 8)),
	1899 => std_logic_vector(to_unsigned(168, 8)),
	1900 => std_logic_vector(to_unsigned(176, 8)),
	1901 => std_logic_vector(to_unsigned(175, 8)),
	1902 => std_logic_vector(to_unsigned(163, 8)),
	1903 => std_logic_vector(to_unsigned(171, 8)),
	1904 => std_logic_vector(to_unsigned(173, 8)),
	1905 => std_logic_vector(to_unsigned(162, 8)),
	1906 => std_logic_vector(to_unsigned(163, 8)),
	1907 => std_logic_vector(to_unsigned(173, 8)),
	1908 => std_logic_vector(to_unsigned(173, 8)),
	1909 => std_logic_vector(to_unsigned(165, 8)),
	1910 => std_logic_vector(to_unsigned(164, 8)),
	1911 => std_logic_vector(to_unsigned(166, 8)),
	1912 => std_logic_vector(to_unsigned(171, 8)),
	1913 => std_logic_vector(to_unsigned(174, 8)),
	1914 => std_logic_vector(to_unsigned(172, 8)),
	1915 => std_logic_vector(to_unsigned(175, 8)),
	1916 => std_logic_vector(to_unsigned(174, 8)),
	1917 => std_logic_vector(to_unsigned(176, 8)),
	1918 => std_logic_vector(to_unsigned(168, 8)),
	1919 => std_logic_vector(to_unsigned(176, 8)),
	1920 => std_logic_vector(to_unsigned(167, 8)),
	1921 => std_logic_vector(to_unsigned(169, 8)),
	1922 => std_logic_vector(to_unsigned(174, 8)),
	1923 => std_logic_vector(to_unsigned(168, 8)),
	1924 => std_logic_vector(to_unsigned(162, 8)),
	1925 => std_logic_vector(to_unsigned(169, 8)),
	1926 => std_logic_vector(to_unsigned(172, 8)),
	1927 => std_logic_vector(to_unsigned(174, 8)),
	1928 => std_logic_vector(to_unsigned(163, 8)),
	1929 => std_logic_vector(to_unsigned(163, 8)),
	1930 => std_logic_vector(to_unsigned(166, 8)),
	1931 => std_logic_vector(to_unsigned(167, 8)),
	1932 => std_logic_vector(to_unsigned(173, 8)),
	1933 => std_logic_vector(to_unsigned(172, 8)),
	1934 => std_logic_vector(to_unsigned(171, 8)),
	1935 => std_logic_vector(to_unsigned(162, 8)),
	1936 => std_logic_vector(to_unsigned(166, 8)),
	1937 => std_logic_vector(to_unsigned(162, 8)),
	1938 => std_logic_vector(to_unsigned(171, 8)),
	1939 => std_logic_vector(to_unsigned(175, 8)),
	1940 => std_logic_vector(to_unsigned(170, 8)),
	1941 => std_logic_vector(to_unsigned(168, 8)),
	1942 => std_logic_vector(to_unsigned(166, 8)),
	1943 => std_logic_vector(to_unsigned(175, 8)),
	1944 => std_logic_vector(to_unsigned(166, 8)),
	1945 => std_logic_vector(to_unsigned(169, 8)),
	1946 => std_logic_vector(to_unsigned(176, 8)),
	1947 => std_logic_vector(to_unsigned(170, 8)),
	1948 => std_logic_vector(to_unsigned(174, 8)),
	1949 => std_logic_vector(to_unsigned(173, 8)),
	1950 => std_logic_vector(to_unsigned(166, 8)),
	1951 => std_logic_vector(to_unsigned(163, 8)),
	1952 => std_logic_vector(to_unsigned(165, 8)),
	1953 => std_logic_vector(to_unsigned(172, 8)),
	1954 => std_logic_vector(to_unsigned(172, 8)),
	1955 => std_logic_vector(to_unsigned(164, 8)),
	1956 => std_logic_vector(to_unsigned(168, 8)),
	1957 => std_logic_vector(to_unsigned(175, 8)),
	1958 => std_logic_vector(to_unsigned(165, 8)),
	1959 => std_logic_vector(to_unsigned(173, 8)),
	1960 => std_logic_vector(to_unsigned(162, 8)),
	1961 => std_logic_vector(to_unsigned(162, 8)),
	1962 => std_logic_vector(to_unsigned(162, 8)),
	1963 => std_logic_vector(to_unsigned(174, 8)),
	1964 => std_logic_vector(to_unsigned(163, 8)),
	1965 => std_logic_vector(to_unsigned(173, 8)),
	1966 => std_logic_vector(to_unsigned(169, 8)),
	1967 => std_logic_vector(to_unsigned(170, 8)),
	1968 => std_logic_vector(to_unsigned(166, 8)),
	1969 => std_logic_vector(to_unsigned(164, 8)),
	1970 => std_logic_vector(to_unsigned(165, 8)),
	1971 => std_logic_vector(to_unsigned(168, 8)),
	1972 => std_logic_vector(to_unsigned(162, 8)),
	1973 => std_logic_vector(to_unsigned(163, 8)),
	1974 => std_logic_vector(to_unsigned(166, 8)),
	1975 => std_logic_vector(to_unsigned(169, 8)),
	1976 => std_logic_vector(to_unsigned(168, 8)),
	1977 => std_logic_vector(to_unsigned(174, 8)),
	1978 => std_logic_vector(to_unsigned(170, 8)),
	1979 => std_logic_vector(to_unsigned(169, 8)),
	1980 => std_logic_vector(to_unsigned(165, 8)),
	1981 => std_logic_vector(to_unsigned(165, 8)),
	1982 => std_logic_vector(to_unsigned(167, 8)),
	1983 => std_logic_vector(to_unsigned(165, 8)),
	1984 => std_logic_vector(to_unsigned(167, 8)),
	1985 => std_logic_vector(to_unsigned(174, 8)),
	1986 => std_logic_vector(to_unsigned(162, 8)),
	1987 => std_logic_vector(to_unsigned(173, 8)),
	1988 => std_logic_vector(to_unsigned(167, 8)),
	1989 => std_logic_vector(to_unsigned(164, 8)),
	1990 => std_logic_vector(to_unsigned(167, 8)),
	1991 => std_logic_vector(to_unsigned(164, 8)),
	1992 => std_logic_vector(to_unsigned(166, 8)),
	1993 => std_logic_vector(to_unsigned(176, 8)),
	1994 => std_logic_vector(to_unsigned(166, 8)),
	1995 => std_logic_vector(to_unsigned(170, 8)),
	1996 => std_logic_vector(to_unsigned(162, 8)),
	1997 => std_logic_vector(to_unsigned(167, 8)),
	1998 => std_logic_vector(to_unsigned(175, 8)),
	1999 => std_logic_vector(to_unsigned(174, 8)),
	2000 => std_logic_vector(to_unsigned(164, 8)),
	2001 => std_logic_vector(to_unsigned(176, 8)),
	2002 => std_logic_vector(to_unsigned(174, 8)),
	2003 => std_logic_vector(to_unsigned(175, 8)),
	2004 => std_logic_vector(to_unsigned(171, 8)),
	2005 => std_logic_vector(to_unsigned(172, 8)),
	2006 => std_logic_vector(to_unsigned(171, 8)),
	2007 => std_logic_vector(to_unsigned(174, 8)),
	2008 => std_logic_vector(to_unsigned(176, 8)),
	2009 => std_logic_vector(to_unsigned(163, 8)),
	2010 => std_logic_vector(to_unsigned(173, 8)),
	2011 => std_logic_vector(to_unsigned(166, 8)),
	2012 => std_logic_vector(to_unsigned(165, 8)),
	2013 => std_logic_vector(to_unsigned(162, 8)),
	2014 => std_logic_vector(to_unsigned(176, 8)),
	2015 => std_logic_vector(to_unsigned(175, 8)),
	2016 => std_logic_vector(to_unsigned(164, 8)),
	2017 => std_logic_vector(to_unsigned(168, 8)),
	2018 => std_logic_vector(to_unsigned(173, 8)),
	2019 => std_logic_vector(to_unsigned(174, 8)),
	2020 => std_logic_vector(to_unsigned(166, 8)),
	2021 => std_logic_vector(to_unsigned(170, 8)),
	2022 => std_logic_vector(to_unsigned(176, 8)),
	2023 => std_logic_vector(to_unsigned(164, 8)),
	2024 => std_logic_vector(to_unsigned(168, 8)),
	2025 => std_logic_vector(to_unsigned(169, 8)),
	2026 => std_logic_vector(to_unsigned(173, 8)),
	2027 => std_logic_vector(to_unsigned(168, 8)),
	2028 => std_logic_vector(to_unsigned(170, 8)),
	2029 => std_logic_vector(to_unsigned(170, 8)),
	2030 => std_logic_vector(to_unsigned(168, 8)),
	2031 => std_logic_vector(to_unsigned(176, 8)),
	2032 => std_logic_vector(to_unsigned(165, 8)),
	2033 => std_logic_vector(to_unsigned(173, 8)),
	2034 => std_logic_vector(to_unsigned(175, 8)),
	2035 => std_logic_vector(to_unsigned(174, 8)),
	2036 => std_logic_vector(to_unsigned(175, 8)),
	2037 => std_logic_vector(to_unsigned(168, 8)),
	2038 => std_logic_vector(to_unsigned(171, 8)),
	2039 => std_logic_vector(to_unsigned(169, 8)),
	2040 => std_logic_vector(to_unsigned(169, 8)),
	2041 => std_logic_vector(to_unsigned(165, 8)),
	2042 => std_logic_vector(to_unsigned(174, 8)),
	2043 => std_logic_vector(to_unsigned(162, 8)),
	2044 => std_logic_vector(to_unsigned(173, 8)),
	2045 => std_logic_vector(to_unsigned(175, 8)),
	2046 => std_logic_vector(to_unsigned(166, 8)),
	2047 => std_logic_vector(to_unsigned(173, 8)),
	2048 => std_logic_vector(to_unsigned(162, 8)),
	2049 => std_logic_vector(to_unsigned(174, 8)),
	2050 => std_logic_vector(to_unsigned(170, 8)),
	2051 => std_logic_vector(to_unsigned(173, 8)),
	2052 => std_logic_vector(to_unsigned(166, 8)),
	2053 => std_logic_vector(to_unsigned(165, 8)),
	2054 => std_logic_vector(to_unsigned(176, 8)),
	2055 => std_logic_vector(to_unsigned(169, 8)),
	2056 => std_logic_vector(to_unsigned(176, 8)),
	2057 => std_logic_vector(to_unsigned(166, 8)),
	2058 => std_logic_vector(to_unsigned(165, 8)),
	2059 => std_logic_vector(to_unsigned(166, 8)),
	2060 => std_logic_vector(to_unsigned(165, 8)),
	2061 => std_logic_vector(to_unsigned(176, 8)),
	2062 => std_logic_vector(to_unsigned(168, 8)),
	2063 => std_logic_vector(to_unsigned(174, 8)),
	2064 => std_logic_vector(to_unsigned(164, 8)),
	2065 => std_logic_vector(to_unsigned(174, 8)),
	2066 => std_logic_vector(to_unsigned(165, 8)),
	2067 => std_logic_vector(to_unsigned(174, 8)),
	2068 => std_logic_vector(to_unsigned(168, 8)),
	2069 => std_logic_vector(to_unsigned(163, 8)),
	2070 => std_logic_vector(to_unsigned(166, 8)),
	2071 => std_logic_vector(to_unsigned(173, 8)),
	2072 => std_logic_vector(to_unsigned(173, 8)),
	2073 => std_logic_vector(to_unsigned(176, 8)),
	2074 => std_logic_vector(to_unsigned(165, 8)),
	2075 => std_logic_vector(to_unsigned(166, 8)),
	2076 => std_logic_vector(to_unsigned(165, 8)),
	2077 => std_logic_vector(to_unsigned(165, 8)),
	2078 => std_logic_vector(to_unsigned(168, 8)),
	2079 => std_logic_vector(to_unsigned(171, 8)),
	2080 => std_logic_vector(to_unsigned(170, 8)),
	2081 => std_logic_vector(to_unsigned(164, 8)),
	2082 => std_logic_vector(to_unsigned(164, 8)),
	2083 => std_logic_vector(to_unsigned(162, 8)),
	2084 => std_logic_vector(to_unsigned(166, 8)),
	2085 => std_logic_vector(to_unsigned(172, 8)),
	2086 => std_logic_vector(to_unsigned(175, 8)),
	2087 => std_logic_vector(to_unsigned(172, 8)),
	2088 => std_logic_vector(to_unsigned(162, 8)),
	2089 => std_logic_vector(to_unsigned(170, 8)),
	2090 => std_logic_vector(to_unsigned(168, 8)),
	2091 => std_logic_vector(to_unsigned(162, 8)),
	2092 => std_logic_vector(to_unsigned(163, 8)),
	2093 => std_logic_vector(to_unsigned(170, 8)),
	2094 => std_logic_vector(to_unsigned(173, 8)),
	2095 => std_logic_vector(to_unsigned(170, 8)),
	2096 => std_logic_vector(to_unsigned(171, 8)),
	2097 => std_logic_vector(to_unsigned(165, 8)),
	2098 => std_logic_vector(to_unsigned(165, 8)),
	2099 => std_logic_vector(to_unsigned(173, 8)),
	2100 => std_logic_vector(to_unsigned(165, 8)),
	2101 => std_logic_vector(to_unsigned(176, 8)),
	2102 => std_logic_vector(to_unsigned(173, 8)),
	2103 => std_logic_vector(to_unsigned(171, 8)),
	2104 => std_logic_vector(to_unsigned(172, 8)),
	2105 => std_logic_vector(to_unsigned(172, 8)),
	2106 => std_logic_vector(to_unsigned(174, 8)),
	2107 => std_logic_vector(to_unsigned(169, 8)),
	2108 => std_logic_vector(to_unsigned(165, 8)),
	2109 => std_logic_vector(to_unsigned(176, 8)),
	2110 => std_logic_vector(to_unsigned(162, 8)),
	2111 => std_logic_vector(to_unsigned(174, 8)),
	2112 => std_logic_vector(to_unsigned(164, 8)),
	2113 => std_logic_vector(to_unsigned(176, 8)),
	2114 => std_logic_vector(to_unsigned(166, 8)),
	2115 => std_logic_vector(to_unsigned(175, 8)),
	2116 => std_logic_vector(to_unsigned(171, 8)),
	2117 => std_logic_vector(to_unsigned(175, 8)),
	2118 => std_logic_vector(to_unsigned(169, 8)),
	2119 => std_logic_vector(to_unsigned(172, 8)),
	2120 => std_logic_vector(to_unsigned(164, 8)),
	2121 => std_logic_vector(to_unsigned(162, 8)),
	2122 => std_logic_vector(to_unsigned(169, 8)),
	2123 => std_logic_vector(to_unsigned(169, 8)),
	2124 => std_logic_vector(to_unsigned(169, 8)),
	2125 => std_logic_vector(to_unsigned(165, 8)),
	2126 => std_logic_vector(to_unsigned(172, 8)),
	2127 => std_logic_vector(to_unsigned(174, 8)),
	2128 => std_logic_vector(to_unsigned(175, 8)),
	2129 => std_logic_vector(to_unsigned(175, 8)),
	2130 => std_logic_vector(to_unsigned(165, 8)),
	2131 => std_logic_vector(to_unsigned(164, 8)),
	2132 => std_logic_vector(to_unsigned(165, 8)),
	2133 => std_logic_vector(to_unsigned(176, 8)),
	2134 => std_logic_vector(to_unsigned(164, 8)),
	2135 => std_logic_vector(to_unsigned(168, 8)),
	2136 => std_logic_vector(to_unsigned(163, 8)),
	2137 => std_logic_vector(to_unsigned(164, 8)),
	2138 => std_logic_vector(to_unsigned(172, 8)),
	2139 => std_logic_vector(to_unsigned(167, 8)),
	2140 => std_logic_vector(to_unsigned(171, 8)),
	2141 => std_logic_vector(to_unsigned(176, 8)),
	2142 => std_logic_vector(to_unsigned(169, 8)),
	2143 => std_logic_vector(to_unsigned(165, 8)),
	2144 => std_logic_vector(to_unsigned(167, 8)),
	2145 => std_logic_vector(to_unsigned(162, 8)),
	2146 => std_logic_vector(to_unsigned(172, 8)),
	2147 => std_logic_vector(to_unsigned(172, 8)),
	2148 => std_logic_vector(to_unsigned(167, 8)),
	2149 => std_logic_vector(to_unsigned(166, 8)),
	2150 => std_logic_vector(to_unsigned(174, 8)),
	2151 => std_logic_vector(to_unsigned(168, 8)),
	2152 => std_logic_vector(to_unsigned(165, 8)),
	2153 => std_logic_vector(to_unsigned(172, 8)),
	2154 => std_logic_vector(to_unsigned(168, 8)),
	2155 => std_logic_vector(to_unsigned(166, 8)),
	2156 => std_logic_vector(to_unsigned(164, 8)),
	2157 => std_logic_vector(to_unsigned(172, 8)),
	2158 => std_logic_vector(to_unsigned(166, 8)),
	2159 => std_logic_vector(to_unsigned(176, 8)),
	2160 => std_logic_vector(to_unsigned(176, 8)),
	2161 => std_logic_vector(to_unsigned(168, 8)),
	2162 => std_logic_vector(to_unsigned(175, 8)),
	2163 => std_logic_vector(to_unsigned(168, 8)),
	2164 => std_logic_vector(to_unsigned(168, 8)),
	2165 => std_logic_vector(to_unsigned(172, 8)),
	2166 => std_logic_vector(to_unsigned(175, 8)),
	2167 => std_logic_vector(to_unsigned(169, 8)),
	2168 => std_logic_vector(to_unsigned(168, 8)),
	2169 => std_logic_vector(to_unsigned(172, 8)),
	2170 => std_logic_vector(to_unsigned(164, 8)),
	2171 => std_logic_vector(to_unsigned(162, 8)),
	2172 => std_logic_vector(to_unsigned(167, 8)),
	2173 => std_logic_vector(to_unsigned(165, 8)),
	2174 => std_logic_vector(to_unsigned(162, 8)),
	2175 => std_logic_vector(to_unsigned(164, 8)),
	2176 => std_logic_vector(to_unsigned(171, 8)),
	2177 => std_logic_vector(to_unsigned(163, 8)),
	2178 => std_logic_vector(to_unsigned(164, 8)),
	2179 => std_logic_vector(to_unsigned(174, 8)),
	2180 => std_logic_vector(to_unsigned(168, 8)),
	2181 => std_logic_vector(to_unsigned(165, 8)),
	2182 => std_logic_vector(to_unsigned(163, 8)),
	2183 => std_logic_vector(to_unsigned(176, 8)),
	2184 => std_logic_vector(to_unsigned(174, 8)),
	2185 => std_logic_vector(to_unsigned(162, 8)),
	2186 => std_logic_vector(to_unsigned(165, 8)),
	2187 => std_logic_vector(to_unsigned(175, 8)),
	2188 => std_logic_vector(to_unsigned(167, 8)),
	2189 => std_logic_vector(to_unsigned(172, 8)),
	2190 => std_logic_vector(to_unsigned(164, 8)),
	2191 => std_logic_vector(to_unsigned(162, 8)),
	2192 => std_logic_vector(to_unsigned(176, 8)),
	2193 => std_logic_vector(to_unsigned(169, 8)),
	2194 => std_logic_vector(to_unsigned(172, 8)),
	2195 => std_logic_vector(to_unsigned(173, 8)),
	2196 => std_logic_vector(to_unsigned(172, 8)),
	2197 => std_logic_vector(to_unsigned(169, 8)),
	2198 => std_logic_vector(to_unsigned(167, 8)),
	2199 => std_logic_vector(to_unsigned(176, 8)),
	2200 => std_logic_vector(to_unsigned(167, 8)),
	2201 => std_logic_vector(to_unsigned(174, 8)),
	2202 => std_logic_vector(to_unsigned(169, 8)),
	2203 => std_logic_vector(to_unsigned(165, 8)),
	2204 => std_logic_vector(to_unsigned(176, 8)),
	2205 => std_logic_vector(to_unsigned(166, 8)),
	2206 => std_logic_vector(to_unsigned(165, 8)),
	2207 => std_logic_vector(to_unsigned(166, 8)),
	2208 => std_logic_vector(to_unsigned(176, 8)),
	2209 => std_logic_vector(to_unsigned(165, 8)),
	2210 => std_logic_vector(to_unsigned(170, 8)),
	2211 => std_logic_vector(to_unsigned(176, 8)),
	2212 => std_logic_vector(to_unsigned(175, 8)),
	2213 => std_logic_vector(to_unsigned(165, 8)),
	2214 => std_logic_vector(to_unsigned(166, 8)),
	2215 => std_logic_vector(to_unsigned(173, 8)),
	2216 => std_logic_vector(to_unsigned(173, 8)),
	2217 => std_logic_vector(to_unsigned(165, 8)),
	2218 => std_logic_vector(to_unsigned(168, 8)),
	2219 => std_logic_vector(to_unsigned(172, 8)),
	2220 => std_logic_vector(to_unsigned(172, 8)),
	2221 => std_logic_vector(to_unsigned(175, 8)),
	2222 => std_logic_vector(to_unsigned(175, 8)),
	2223 => std_logic_vector(to_unsigned(162, 8)),
	2224 => std_logic_vector(to_unsigned(163, 8)),
	2225 => std_logic_vector(to_unsigned(165, 8)),
	2226 => std_logic_vector(to_unsigned(174, 8)),
	2227 => std_logic_vector(to_unsigned(167, 8)),
	2228 => std_logic_vector(to_unsigned(173, 8)),
	2229 => std_logic_vector(to_unsigned(176, 8)),
	2230 => std_logic_vector(to_unsigned(173, 8)),
	2231 => std_logic_vector(to_unsigned(163, 8)),
	2232 => std_logic_vector(to_unsigned(175, 8)),
	2233 => std_logic_vector(to_unsigned(175, 8)),
	2234 => std_logic_vector(to_unsigned(168, 8)),
	2235 => std_logic_vector(to_unsigned(168, 8)),
	2236 => std_logic_vector(to_unsigned(164, 8)),
	2237 => std_logic_vector(to_unsigned(164, 8)),
	2238 => std_logic_vector(to_unsigned(170, 8)),
	2239 => std_logic_vector(to_unsigned(174, 8)),
	2240 => std_logic_vector(to_unsigned(168, 8)),
	2241 => std_logic_vector(to_unsigned(175, 8)),
	2242 => std_logic_vector(to_unsigned(166, 8)),
	2243 => std_logic_vector(to_unsigned(174, 8)),
	2244 => std_logic_vector(to_unsigned(162, 8)),
	2245 => std_logic_vector(to_unsigned(167, 8)),
	2246 => std_logic_vector(to_unsigned(164, 8)),
	2247 => std_logic_vector(to_unsigned(168, 8)),
	2248 => std_logic_vector(to_unsigned(169, 8)),
	2249 => std_logic_vector(to_unsigned(176, 8)),
	2250 => std_logic_vector(to_unsigned(172, 8)),
	2251 => std_logic_vector(to_unsigned(169, 8)),
	2252 => std_logic_vector(to_unsigned(166, 8)),
	2253 => std_logic_vector(to_unsigned(169, 8)),
	2254 => std_logic_vector(to_unsigned(176, 8)),
	2255 => std_logic_vector(to_unsigned(162, 8)),
	2256 => std_logic_vector(to_unsigned(164, 8)),
	2257 => std_logic_vector(to_unsigned(172, 8)),
	2258 => std_logic_vector(to_unsigned(176, 8)),
	2259 => std_logic_vector(to_unsigned(166, 8)),
	2260 => std_logic_vector(to_unsigned(169, 8)),
	2261 => std_logic_vector(to_unsigned(167, 8)),
	2262 => std_logic_vector(to_unsigned(165, 8)),
	2263 => std_logic_vector(to_unsigned(162, 8)),
	2264 => std_logic_vector(to_unsigned(176, 8)),
	2265 => std_logic_vector(to_unsigned(164, 8)),
	2266 => std_logic_vector(to_unsigned(172, 8)),
	2267 => std_logic_vector(to_unsigned(175, 8)),
	2268 => std_logic_vector(to_unsigned(164, 8)),
	2269 => std_logic_vector(to_unsigned(163, 8)),
	2270 => std_logic_vector(to_unsigned(165, 8)),
	2271 => std_logic_vector(to_unsigned(165, 8)),
	2272 => std_logic_vector(to_unsigned(167, 8)),
	2273 => std_logic_vector(to_unsigned(173, 8)),
	2274 => std_logic_vector(to_unsigned(170, 8)),
	2275 => std_logic_vector(to_unsigned(175, 8)),
	2276 => std_logic_vector(to_unsigned(172, 8)),
	2277 => std_logic_vector(to_unsigned(165, 8)),
	2278 => std_logic_vector(to_unsigned(165, 8)),
	2279 => std_logic_vector(to_unsigned(175, 8)),
	2280 => std_logic_vector(to_unsigned(176, 8)),
	2281 => std_logic_vector(to_unsigned(169, 8)),
	2282 => std_logic_vector(to_unsigned(162, 8)),
	2283 => std_logic_vector(to_unsigned(173, 8)),
	2284 => std_logic_vector(to_unsigned(167, 8)),
	2285 => std_logic_vector(to_unsigned(172, 8)),
	2286 => std_logic_vector(to_unsigned(174, 8)),
	2287 => std_logic_vector(to_unsigned(166, 8)),
	2288 => std_logic_vector(to_unsigned(165, 8)),
	2289 => std_logic_vector(to_unsigned(169, 8)),
	2290 => std_logic_vector(to_unsigned(169, 8)),
	2291 => std_logic_vector(to_unsigned(169, 8)),
	2292 => std_logic_vector(to_unsigned(171, 8)),
	2293 => std_logic_vector(to_unsigned(173, 8)),
	2294 => std_logic_vector(to_unsigned(174, 8)),
	2295 => std_logic_vector(to_unsigned(164, 8)),
	2296 => std_logic_vector(to_unsigned(168, 8)),
	2297 => std_logic_vector(to_unsigned(175, 8)),
	2298 => std_logic_vector(to_unsigned(174, 8)),
	2299 => std_logic_vector(to_unsigned(174, 8)),
	2300 => std_logic_vector(to_unsigned(164, 8)),
	2301 => std_logic_vector(to_unsigned(170, 8)),
	2302 => std_logic_vector(to_unsigned(163, 8)),
	2303 => std_logic_vector(to_unsigned(174, 8)),
	2304 => std_logic_vector(to_unsigned(168, 8)),
	2305 => std_logic_vector(to_unsigned(166, 8)),
	2306 => std_logic_vector(to_unsigned(162, 8)),
	2307 => std_logic_vector(to_unsigned(176, 8)),
	2308 => std_logic_vector(to_unsigned(170, 8)),
	2309 => std_logic_vector(to_unsigned(166, 8)),
	2310 => std_logic_vector(to_unsigned(173, 8)),
	2311 => std_logic_vector(to_unsigned(168, 8)),
	2312 => std_logic_vector(to_unsigned(173, 8)),
	2313 => std_logic_vector(to_unsigned(175, 8)),
	2314 => std_logic_vector(to_unsigned(166, 8)),
	2315 => std_logic_vector(to_unsigned(168, 8)),
	2316 => std_logic_vector(to_unsigned(168, 8)),
	2317 => std_logic_vector(to_unsigned(170, 8)),
	2318 => std_logic_vector(to_unsigned(164, 8)),
	2319 => std_logic_vector(to_unsigned(162, 8)),
	2320 => std_logic_vector(to_unsigned(168, 8)),
	2321 => std_logic_vector(to_unsigned(164, 8)),
	2322 => std_logic_vector(to_unsigned(173, 8)),
	2323 => std_logic_vector(to_unsigned(163, 8)),
	2324 => std_logic_vector(to_unsigned(170, 8)),
	2325 => std_logic_vector(to_unsigned(166, 8)),
	2326 => std_logic_vector(to_unsigned(173, 8)),
	2327 => std_logic_vector(to_unsigned(170, 8)),
	2328 => std_logic_vector(to_unsigned(169, 8)),
	2329 => std_logic_vector(to_unsigned(162, 8)),
	2330 => std_logic_vector(to_unsigned(172, 8)),
	2331 => std_logic_vector(to_unsigned(174, 8)),
	2332 => std_logic_vector(to_unsigned(164, 8)),
	2333 => std_logic_vector(to_unsigned(166, 8)),
	2334 => std_logic_vector(to_unsigned(171, 8)),
	2335 => std_logic_vector(to_unsigned(171, 8)),
	2336 => std_logic_vector(to_unsigned(174, 8)),
	2337 => std_logic_vector(to_unsigned(164, 8)),
	2338 => std_logic_vector(to_unsigned(174, 8)),
	2339 => std_logic_vector(to_unsigned(175, 8)),
	2340 => std_logic_vector(to_unsigned(167, 8)),
	2341 => std_logic_vector(to_unsigned(176, 8)),
	2342 => std_logic_vector(to_unsigned(172, 8)),
	2343 => std_logic_vector(to_unsigned(163, 8)),
	2344 => std_logic_vector(to_unsigned(174, 8)),
	2345 => std_logic_vector(to_unsigned(175, 8)),
	2346 => std_logic_vector(to_unsigned(162, 8)),
	2347 => std_logic_vector(to_unsigned(173, 8)),
	2348 => std_logic_vector(to_unsigned(172, 8)),
	2349 => std_logic_vector(to_unsigned(166, 8)),
	2350 => std_logic_vector(to_unsigned(170, 8)),
	2351 => std_logic_vector(to_unsigned(171, 8)),
	2352 => std_logic_vector(to_unsigned(163, 8)),
	2353 => std_logic_vector(to_unsigned(162, 8)),
	2354 => std_logic_vector(to_unsigned(169, 8)),
	2355 => std_logic_vector(to_unsigned(176, 8)),
	2356 => std_logic_vector(to_unsigned(170, 8)),
	2357 => std_logic_vector(to_unsigned(162, 8)),
	2358 => std_logic_vector(to_unsigned(169, 8)),
	2359 => std_logic_vector(to_unsigned(173, 8)),
	2360 => std_logic_vector(to_unsigned(173, 8)),
	2361 => std_logic_vector(to_unsigned(170, 8)),
	2362 => std_logic_vector(to_unsigned(170, 8)),
	2363 => std_logic_vector(to_unsigned(165, 8)),
	2364 => std_logic_vector(to_unsigned(175, 8)),
	2365 => std_logic_vector(to_unsigned(162, 8)),
	2366 => std_logic_vector(to_unsigned(171, 8)),
	2367 => std_logic_vector(to_unsigned(164, 8)),
	2368 => std_logic_vector(to_unsigned(162, 8)),
	2369 => std_logic_vector(to_unsigned(170, 8)),
	2370 => std_logic_vector(to_unsigned(162, 8)),
	2371 => std_logic_vector(to_unsigned(166, 8)),
	2372 => std_logic_vector(to_unsigned(176, 8)),
	2373 => std_logic_vector(to_unsigned(165, 8)),
	2374 => std_logic_vector(to_unsigned(172, 8)),
	2375 => std_logic_vector(to_unsigned(167, 8)),
	2376 => std_logic_vector(to_unsigned(173, 8)),
	2377 => std_logic_vector(to_unsigned(165, 8)),
	2378 => std_logic_vector(to_unsigned(162, 8)),
	2379 => std_logic_vector(to_unsigned(174, 8)),
	2380 => std_logic_vector(to_unsigned(173, 8)),
	2381 => std_logic_vector(to_unsigned(162, 8)),
	2382 => std_logic_vector(to_unsigned(166, 8)),
	2383 => std_logic_vector(to_unsigned(165, 8)),
	2384 => std_logic_vector(to_unsigned(168, 8)),
	2385 => std_logic_vector(to_unsigned(163, 8)),
	2386 => std_logic_vector(to_unsigned(165, 8)),
	2387 => std_logic_vector(to_unsigned(163, 8)),
	2388 => std_logic_vector(to_unsigned(170, 8)),
	2389 => std_logic_vector(to_unsigned(163, 8)),
	2390 => std_logic_vector(to_unsigned(167, 8)),
	2391 => std_logic_vector(to_unsigned(169, 8)),
	2392 => std_logic_vector(to_unsigned(175, 8)),
	2393 => std_logic_vector(to_unsigned(164, 8)),
	2394 => std_logic_vector(to_unsigned(164, 8)),
	2395 => std_logic_vector(to_unsigned(168, 8)),
	2396 => std_logic_vector(to_unsigned(176, 8)),
	2397 => std_logic_vector(to_unsigned(162, 8)),
	2398 => std_logic_vector(to_unsigned(163, 8)),
	2399 => std_logic_vector(to_unsigned(169, 8)),
	2400 => std_logic_vector(to_unsigned(162, 8)),
	2401 => std_logic_vector(to_unsigned(166, 8)),
	2402 => std_logic_vector(to_unsigned(162, 8)),
	2403 => std_logic_vector(to_unsigned(164, 8)),
	2404 => std_logic_vector(to_unsigned(169, 8)),
	2405 => std_logic_vector(to_unsigned(162, 8)),
	2406 => std_logic_vector(to_unsigned(166, 8)),
	2407 => std_logic_vector(to_unsigned(175, 8)),
	2408 => std_logic_vector(to_unsigned(175, 8)),
	2409 => std_logic_vector(to_unsigned(166, 8)),
	2410 => std_logic_vector(to_unsigned(167, 8)),
	2411 => std_logic_vector(to_unsigned(172, 8)),
	2412 => std_logic_vector(to_unsigned(166, 8)),
	2413 => std_logic_vector(to_unsigned(172, 8)),
	2414 => std_logic_vector(to_unsigned(169, 8)),
	2415 => std_logic_vector(to_unsigned(176, 8)),
	2416 => std_logic_vector(to_unsigned(163, 8)),
	2417 => std_logic_vector(to_unsigned(175, 8)),
	2418 => std_logic_vector(to_unsigned(163, 8)),
	2419 => std_logic_vector(to_unsigned(169, 8)),
	2420 => std_logic_vector(to_unsigned(166, 8)),
	2421 => std_logic_vector(to_unsigned(164, 8)),
	2422 => std_logic_vector(to_unsigned(170, 8)),
	2423 => std_logic_vector(to_unsigned(164, 8)),
	2424 => std_logic_vector(to_unsigned(171, 8)),
	2425 => std_logic_vector(to_unsigned(174, 8)),
	2426 => std_logic_vector(to_unsigned(173, 8)),
	2427 => std_logic_vector(to_unsigned(163, 8)),
	2428 => std_logic_vector(to_unsigned(162, 8)),
	2429 => std_logic_vector(to_unsigned(175, 8)),
	2430 => std_logic_vector(to_unsigned(163, 8)),
	2431 => std_logic_vector(to_unsigned(173, 8)),
	2432 => std_logic_vector(to_unsigned(174, 8)),
	2433 => std_logic_vector(to_unsigned(165, 8)),
	2434 => std_logic_vector(to_unsigned(164, 8)),
	2435 => std_logic_vector(to_unsigned(174, 8)),
	2436 => std_logic_vector(to_unsigned(165, 8)),
	2437 => std_logic_vector(to_unsigned(162, 8)),
	2438 => std_logic_vector(to_unsigned(167, 8)),
	2439 => std_logic_vector(to_unsigned(170, 8)),
	2440 => std_logic_vector(to_unsigned(163, 8)),
	2441 => std_logic_vector(to_unsigned(173, 8)),
	2442 => std_logic_vector(to_unsigned(171, 8)),
	2443 => std_logic_vector(to_unsigned(174, 8)),
	2444 => std_logic_vector(to_unsigned(173, 8)),
	2445 => std_logic_vector(to_unsigned(165, 8)),
	2446 => std_logic_vector(to_unsigned(170, 8)),
	2447 => std_logic_vector(to_unsigned(174, 8)),
	2448 => std_logic_vector(to_unsigned(172, 8)),
	2449 => std_logic_vector(to_unsigned(176, 8)),
	2450 => std_logic_vector(to_unsigned(175, 8)),
	2451 => std_logic_vector(to_unsigned(167, 8)),
	2452 => std_logic_vector(to_unsigned(166, 8)),
	2453 => std_logic_vector(to_unsigned(172, 8)),
	2454 => std_logic_vector(to_unsigned(166, 8)),
	2455 => std_logic_vector(to_unsigned(165, 8)),
	2456 => std_logic_vector(to_unsigned(167, 8)),
	2457 => std_logic_vector(to_unsigned(168, 8)),
	2458 => std_logic_vector(to_unsigned(173, 8)),
	2459 => std_logic_vector(to_unsigned(164, 8)),
	2460 => std_logic_vector(to_unsigned(167, 8)),
	2461 => std_logic_vector(to_unsigned(163, 8)),
	2462 => std_logic_vector(to_unsigned(166, 8)),
	2463 => std_logic_vector(to_unsigned(174, 8)),
	2464 => std_logic_vector(to_unsigned(174, 8)),
	2465 => std_logic_vector(to_unsigned(164, 8)),
	2466 => std_logic_vector(to_unsigned(171, 8)),
	2467 => std_logic_vector(to_unsigned(168, 8)),
	2468 => std_logic_vector(to_unsigned(165, 8)),
	2469 => std_logic_vector(to_unsigned(168, 8)),
	2470 => std_logic_vector(to_unsigned(175, 8)),
	2471 => std_logic_vector(to_unsigned(174, 8)),
	2472 => std_logic_vector(to_unsigned(174, 8)),
	2473 => std_logic_vector(to_unsigned(165, 8)),
	2474 => std_logic_vector(to_unsigned(163, 8)),
	2475 => std_logic_vector(to_unsigned(176, 8)),
	2476 => std_logic_vector(to_unsigned(169, 8)),
	2477 => std_logic_vector(to_unsigned(172, 8)),
	2478 => std_logic_vector(to_unsigned(171, 8)),
	2479 => std_logic_vector(to_unsigned(163, 8)),
	2480 => std_logic_vector(to_unsigned(171, 8)),
	2481 => std_logic_vector(to_unsigned(165, 8)),
	2482 => std_logic_vector(to_unsigned(173, 8)),
	2483 => std_logic_vector(to_unsigned(166, 8)),
	2484 => std_logic_vector(to_unsigned(171, 8)),
	2485 => std_logic_vector(to_unsigned(173, 8)),
	2486 => std_logic_vector(to_unsigned(164, 8)),
	2487 => std_logic_vector(to_unsigned(169, 8)),
	2488 => std_logic_vector(to_unsigned(163, 8)),
	2489 => std_logic_vector(to_unsigned(175, 8)),
	2490 => std_logic_vector(to_unsigned(172, 8)),
	2491 => std_logic_vector(to_unsigned(166, 8)),
	2492 => std_logic_vector(to_unsigned(175, 8)),
	2493 => std_logic_vector(to_unsigned(167, 8)),
	2494 => std_logic_vector(to_unsigned(173, 8)),
	2495 => std_logic_vector(to_unsigned(164, 8)),
	2496 => std_logic_vector(to_unsigned(166, 8)),
	2497 => std_logic_vector(to_unsigned(169, 8)),
	2498 => std_logic_vector(to_unsigned(172, 8)),
	2499 => std_logic_vector(to_unsigned(169, 8)),
	2500 => std_logic_vector(to_unsigned(175, 8)),
	2501 => std_logic_vector(to_unsigned(162, 8)),
	2502 => std_logic_vector(to_unsigned(175, 8)),
	2503 => std_logic_vector(to_unsigned(167, 8)),
	2504 => std_logic_vector(to_unsigned(175, 8)),
	2505 => std_logic_vector(to_unsigned(170, 8)),
	2506 => std_logic_vector(to_unsigned(175, 8)),
	2507 => std_logic_vector(to_unsigned(175, 8)),
	2508 => std_logic_vector(to_unsigned(176, 8)),
	2509 => std_logic_vector(to_unsigned(169, 8)),
	2510 => std_logic_vector(to_unsigned(174, 8)),
	2511 => std_logic_vector(to_unsigned(172, 8)),
	2512 => std_logic_vector(to_unsigned(162, 8)),
	2513 => std_logic_vector(to_unsigned(162, 8)),
	2514 => std_logic_vector(to_unsigned(172, 8)),
	2515 => std_logic_vector(to_unsigned(174, 8)),
	2516 => std_logic_vector(to_unsigned(167, 8)),
	2517 => std_logic_vector(to_unsigned(164, 8)),
	2518 => std_logic_vector(to_unsigned(175, 8)),
	2519 => std_logic_vector(to_unsigned(174, 8)),
	2520 => std_logic_vector(to_unsigned(173, 8)),
	2521 => std_logic_vector(to_unsigned(167, 8)),
	2522 => std_logic_vector(to_unsigned(164, 8)),
	2523 => std_logic_vector(to_unsigned(172, 8)),
	2524 => std_logic_vector(to_unsigned(168, 8)),
	2525 => std_logic_vector(to_unsigned(170, 8)),
	2526 => std_logic_vector(to_unsigned(176, 8)),
	2527 => std_logic_vector(to_unsigned(175, 8)),
	2528 => std_logic_vector(to_unsigned(163, 8)),
	2529 => std_logic_vector(to_unsigned(163, 8)),
	2530 => std_logic_vector(to_unsigned(168, 8)),
	2531 => std_logic_vector(to_unsigned(169, 8)),
	2532 => std_logic_vector(to_unsigned(172, 8)),
	2533 => std_logic_vector(to_unsigned(176, 8)),
	2534 => std_logic_vector(to_unsigned(163, 8)),
	2535 => std_logic_vector(to_unsigned(174, 8)),
	2536 => std_logic_vector(to_unsigned(174, 8)),
	2537 => std_logic_vector(to_unsigned(169, 8)),
	2538 => std_logic_vector(to_unsigned(175, 8)),
	2539 => std_logic_vector(to_unsigned(173, 8)),
	2540 => std_logic_vector(to_unsigned(173, 8)),
	2541 => std_logic_vector(to_unsigned(169, 8)),
	2542 => std_logic_vector(to_unsigned(170, 8)),
	2543 => std_logic_vector(to_unsigned(169, 8)),
	2544 => std_logic_vector(to_unsigned(172, 8)),
	2545 => std_logic_vector(to_unsigned(172, 8)),
	2546 => std_logic_vector(to_unsigned(166, 8)),
	2547 => std_logic_vector(to_unsigned(171, 8)),
	2548 => std_logic_vector(to_unsigned(167, 8)),
	2549 => std_logic_vector(to_unsigned(172, 8)),
	2550 => std_logic_vector(to_unsigned(173, 8)),
	2551 => std_logic_vector(to_unsigned(175, 8)),
	2552 => std_logic_vector(to_unsigned(169, 8)),
	2553 => std_logic_vector(to_unsigned(165, 8)),
	2554 => std_logic_vector(to_unsigned(172, 8)),
	2555 => std_logic_vector(to_unsigned(165, 8)),
	2556 => std_logic_vector(to_unsigned(169, 8)),
	2557 => std_logic_vector(to_unsigned(163, 8)),
	2558 => std_logic_vector(to_unsigned(168, 8)),
	2559 => std_logic_vector(to_unsigned(165, 8)),
	2560 => std_logic_vector(to_unsigned(162, 8)),
	2561 => std_logic_vector(to_unsigned(168, 8)),
	2562 => std_logic_vector(to_unsigned(174, 8)),
	2563 => std_logic_vector(to_unsigned(175, 8)),
	2564 => std_logic_vector(to_unsigned(168, 8)),
	2565 => std_logic_vector(to_unsigned(164, 8)),
	2566 => std_logic_vector(to_unsigned(168, 8)),
	2567 => std_logic_vector(to_unsigned(166, 8)),
	2568 => std_logic_vector(to_unsigned(176, 8)),
	2569 => std_logic_vector(to_unsigned(173, 8)),
	2570 => std_logic_vector(to_unsigned(172, 8)),
	2571 => std_logic_vector(to_unsigned(173, 8)),
	2572 => std_logic_vector(to_unsigned(168, 8)),
	2573 => std_logic_vector(to_unsigned(172, 8)),
	2574 => std_logic_vector(to_unsigned(173, 8)),
	2575 => std_logic_vector(to_unsigned(172, 8)),
	2576 => std_logic_vector(to_unsigned(171, 8)),
	2577 => std_logic_vector(to_unsigned(176, 8)),
	2578 => std_logic_vector(to_unsigned(167, 8)),
	2579 => std_logic_vector(to_unsigned(174, 8)),
	2580 => std_logic_vector(to_unsigned(164, 8)),
	2581 => std_logic_vector(to_unsigned(162, 8)),
	2582 => std_logic_vector(to_unsigned(172, 8)),
	2583 => std_logic_vector(to_unsigned(172, 8)),
	2584 => std_logic_vector(to_unsigned(169, 8)),
	2585 => std_logic_vector(to_unsigned(162, 8)),
	2586 => std_logic_vector(to_unsigned(165, 8)),
	2587 => std_logic_vector(to_unsigned(175, 8)),
	2588 => std_logic_vector(to_unsigned(169, 8)),
	2589 => std_logic_vector(to_unsigned(168, 8)),
	2590 => std_logic_vector(to_unsigned(169, 8)),
	2591 => std_logic_vector(to_unsigned(172, 8)),
	2592 => std_logic_vector(to_unsigned(163, 8)),
	2593 => std_logic_vector(to_unsigned(165, 8)),
	2594 => std_logic_vector(to_unsigned(164, 8)),
	2595 => std_logic_vector(to_unsigned(174, 8)),
	2596 => std_logic_vector(to_unsigned(166, 8)),
	2597 => std_logic_vector(to_unsigned(164, 8)),
	2598 => std_logic_vector(to_unsigned(176, 8)),
	2599 => std_logic_vector(to_unsigned(172, 8)),
	2600 => std_logic_vector(to_unsigned(166, 8)),
	2601 => std_logic_vector(to_unsigned(164, 8)),
	2602 => std_logic_vector(to_unsigned(162, 8)),
	2603 => std_logic_vector(to_unsigned(165, 8)),
	2604 => std_logic_vector(to_unsigned(165, 8)),
	2605 => std_logic_vector(to_unsigned(167, 8)),
	2606 => std_logic_vector(to_unsigned(167, 8)),
	2607 => std_logic_vector(to_unsigned(174, 8)),
	2608 => std_logic_vector(to_unsigned(165, 8)),
	2609 => std_logic_vector(to_unsigned(172, 8)),
	2610 => std_logic_vector(to_unsigned(165, 8)),
	2611 => std_logic_vector(to_unsigned(167, 8)),
	2612 => std_logic_vector(to_unsigned(164, 8)),
	2613 => std_logic_vector(to_unsigned(174, 8)),
	2614 => std_logic_vector(to_unsigned(164, 8)),
	2615 => std_logic_vector(to_unsigned(166, 8)),
	2616 => std_logic_vector(to_unsigned(170, 8)),
	2617 => std_logic_vector(to_unsigned(173, 8)),
	2618 => std_logic_vector(to_unsigned(168, 8)),
	2619 => std_logic_vector(to_unsigned(173, 8)),
	2620 => std_logic_vector(to_unsigned(164, 8)),
	2621 => std_logic_vector(to_unsigned(164, 8)),
	2622 => std_logic_vector(to_unsigned(165, 8)),
	2623 => std_logic_vector(to_unsigned(170, 8)),
	2624 => std_logic_vector(to_unsigned(171, 8)),
	2625 => std_logic_vector(to_unsigned(164, 8)),
	2626 => std_logic_vector(to_unsigned(162, 8)),
	2627 => std_logic_vector(to_unsigned(166, 8)),
	2628 => std_logic_vector(to_unsigned(174, 8)),
	2629 => std_logic_vector(to_unsigned(167, 8)),
	2630 => std_logic_vector(to_unsigned(166, 8)),
	2631 => std_logic_vector(to_unsigned(166, 8)),
	2632 => std_logic_vector(to_unsigned(170, 8)),
	2633 => std_logic_vector(to_unsigned(171, 8)),
	2634 => std_logic_vector(to_unsigned(164, 8)),
	2635 => std_logic_vector(to_unsigned(169, 8)),
	2636 => std_logic_vector(to_unsigned(171, 8)),
	2637 => std_logic_vector(to_unsigned(169, 8)),
	2638 => std_logic_vector(to_unsigned(164, 8)),
	2639 => std_logic_vector(to_unsigned(172, 8)),
	2640 => std_logic_vector(to_unsigned(171, 8)),
	2641 => std_logic_vector(to_unsigned(173, 8)),
	2642 => std_logic_vector(to_unsigned(172, 8)),
	2643 => std_logic_vector(to_unsigned(173, 8)),
	2644 => std_logic_vector(to_unsigned(164, 8)),
	2645 => std_logic_vector(to_unsigned(170, 8)),
	2646 => std_logic_vector(to_unsigned(170, 8)),
	2647 => std_logic_vector(to_unsigned(167, 8)),
	2648 => std_logic_vector(to_unsigned(167, 8)),
	2649 => std_logic_vector(to_unsigned(173, 8)),
	2650 => std_logic_vector(to_unsigned(162, 8)),
	2651 => std_logic_vector(to_unsigned(176, 8)),
	2652 => std_logic_vector(to_unsigned(165, 8)),
	2653 => std_logic_vector(to_unsigned(162, 8)),
	2654 => std_logic_vector(to_unsigned(163, 8)),
	2655 => std_logic_vector(to_unsigned(162, 8)),
	2656 => std_logic_vector(to_unsigned(163, 8)),
	2657 => std_logic_vector(to_unsigned(169, 8)),
	2658 => std_logic_vector(to_unsigned(172, 8)),
	2659 => std_logic_vector(to_unsigned(175, 8)),
	2660 => std_logic_vector(to_unsigned(168, 8)),
	2661 => std_logic_vector(to_unsigned(176, 8)),
	2662 => std_logic_vector(to_unsigned(173, 8)),
	2663 => std_logic_vector(to_unsigned(175, 8)),
	2664 => std_logic_vector(to_unsigned(168, 8)),
	2665 => std_logic_vector(to_unsigned(165, 8)),
	2666 => std_logic_vector(to_unsigned(169, 8)),
	2667 => std_logic_vector(to_unsigned(164, 8)),
	2668 => std_logic_vector(to_unsigned(163, 8)),
	2669 => std_logic_vector(to_unsigned(162, 8)),
	2670 => std_logic_vector(to_unsigned(167, 8)),
	2671 => std_logic_vector(to_unsigned(166, 8)),
	2672 => std_logic_vector(to_unsigned(173, 8)),
	2673 => std_logic_vector(to_unsigned(169, 8)),
	2674 => std_logic_vector(to_unsigned(169, 8)),
	2675 => std_logic_vector(to_unsigned(166, 8)),
	2676 => std_logic_vector(to_unsigned(167, 8)),
	2677 => std_logic_vector(to_unsigned(171, 8)),
	2678 => std_logic_vector(to_unsigned(175, 8)),
	2679 => std_logic_vector(to_unsigned(166, 8)),
	2680 => std_logic_vector(to_unsigned(172, 8)),
	2681 => std_logic_vector(to_unsigned(172, 8)),
	2682 => std_logic_vector(to_unsigned(172, 8)),
	2683 => std_logic_vector(to_unsigned(175, 8)),
	2684 => std_logic_vector(to_unsigned(176, 8)),
	2685 => std_logic_vector(to_unsigned(166, 8)),
	2686 => std_logic_vector(to_unsigned(175, 8)),
	2687 => std_logic_vector(to_unsigned(169, 8)),
	2688 => std_logic_vector(to_unsigned(165, 8)),
	2689 => std_logic_vector(to_unsigned(176, 8)),
	2690 => std_logic_vector(to_unsigned(170, 8)),
	2691 => std_logic_vector(to_unsigned(172, 8)),
	2692 => std_logic_vector(to_unsigned(173, 8)),
	2693 => std_logic_vector(to_unsigned(166, 8)),
	2694 => std_logic_vector(to_unsigned(163, 8)),
	2695 => std_logic_vector(to_unsigned(166, 8)),
	2696 => std_logic_vector(to_unsigned(165, 8)),
	2697 => std_logic_vector(to_unsigned(175, 8)),
	2698 => std_logic_vector(to_unsigned(168, 8)),
	2699 => std_logic_vector(to_unsigned(174, 8)),
	2700 => std_logic_vector(to_unsigned(167, 8)),
	2701 => std_logic_vector(to_unsigned(174, 8)),
	2702 => std_logic_vector(to_unsigned(169, 8)),
	2703 => std_logic_vector(to_unsigned(173, 8)),
	2704 => std_logic_vector(to_unsigned(169, 8)),
	2705 => std_logic_vector(to_unsigned(163, 8)),
	2706 => std_logic_vector(to_unsigned(168, 8)),
	2707 => std_logic_vector(to_unsigned(168, 8)),
	2708 => std_logic_vector(to_unsigned(162, 8)),
	2709 => std_logic_vector(to_unsigned(171, 8)),
	2710 => std_logic_vector(to_unsigned(168, 8)),
	2711 => std_logic_vector(to_unsigned(163, 8)),
	2712 => std_logic_vector(to_unsigned(176, 8)),
	2713 => std_logic_vector(to_unsigned(174, 8)),
	2714 => std_logic_vector(to_unsigned(169, 8)),
	2715 => std_logic_vector(to_unsigned(175, 8)),
	2716 => std_logic_vector(to_unsigned(169, 8)),
	2717 => std_logic_vector(to_unsigned(164, 8)),
	2718 => std_logic_vector(to_unsigned(175, 8)),
	2719 => std_logic_vector(to_unsigned(172, 8)),
	2720 => std_logic_vector(to_unsigned(170, 8)),
	2721 => std_logic_vector(to_unsigned(166, 8)),
	2722 => std_logic_vector(to_unsigned(175, 8)),
	2723 => std_logic_vector(to_unsigned(164, 8)),
	2724 => std_logic_vector(to_unsigned(167, 8)),
	2725 => std_logic_vector(to_unsigned(173, 8)),
	2726 => std_logic_vector(to_unsigned(172, 8)),
	2727 => std_logic_vector(to_unsigned(171, 8)),
	2728 => std_logic_vector(to_unsigned(175, 8)),
	2729 => std_logic_vector(to_unsigned(172, 8)),
	2730 => std_logic_vector(to_unsigned(166, 8)),
	2731 => std_logic_vector(to_unsigned(162, 8)),
	2732 => std_logic_vector(to_unsigned(166, 8)),
	2733 => std_logic_vector(to_unsigned(166, 8)),
	2734 => std_logic_vector(to_unsigned(165, 8)),
	2735 => std_logic_vector(to_unsigned(171, 8)),
	2736 => std_logic_vector(to_unsigned(167, 8)),
	2737 => std_logic_vector(to_unsigned(176, 8)),
	2738 => std_logic_vector(to_unsigned(175, 8)),
	2739 => std_logic_vector(to_unsigned(173, 8)),
	2740 => std_logic_vector(to_unsigned(167, 8)),
	2741 => std_logic_vector(to_unsigned(165, 8)),
	2742 => std_logic_vector(to_unsigned(165, 8)),
	2743 => std_logic_vector(to_unsigned(168, 8)),
	2744 => std_logic_vector(to_unsigned(166, 8)),
	2745 => std_logic_vector(to_unsigned(164, 8)),
	2746 => std_logic_vector(to_unsigned(171, 8)),
	2747 => std_logic_vector(to_unsigned(175, 8)),
	2748 => std_logic_vector(to_unsigned(168, 8)),
	2749 => std_logic_vector(to_unsigned(176, 8)),
	2750 => std_logic_vector(to_unsigned(171, 8)),
	2751 => std_logic_vector(to_unsigned(169, 8)),
	2752 => std_logic_vector(to_unsigned(167, 8)),
	2753 => std_logic_vector(to_unsigned(167, 8)),
	2754 => std_logic_vector(to_unsigned(174, 8)),
	2755 => std_logic_vector(to_unsigned(167, 8)),
	2756 => std_logic_vector(to_unsigned(174, 8)),
	2757 => std_logic_vector(to_unsigned(167, 8)),
	2758 => std_logic_vector(to_unsigned(172, 8)),
	2759 => std_logic_vector(to_unsigned(171, 8)),
	2760 => std_logic_vector(to_unsigned(165, 8)),
	2761 => std_logic_vector(to_unsigned(171, 8)),
	2762 => std_logic_vector(to_unsigned(176, 8)),
	2763 => std_logic_vector(to_unsigned(170, 8)),
	2764 => std_logic_vector(to_unsigned(163, 8)),
	2765 => std_logic_vector(to_unsigned(172, 8)),
	2766 => std_logic_vector(to_unsigned(172, 8)),
	2767 => std_logic_vector(to_unsigned(170, 8)),
	2768 => std_logic_vector(to_unsigned(168, 8)),
	2769 => std_logic_vector(to_unsigned(168, 8)),
	2770 => std_logic_vector(to_unsigned(171, 8)),
	2771 => std_logic_vector(to_unsigned(173, 8)),
	2772 => std_logic_vector(to_unsigned(172, 8)),
	2773 => std_logic_vector(to_unsigned(168, 8)),
	2774 => std_logic_vector(to_unsigned(175, 8)),
	2775 => std_logic_vector(to_unsigned(165, 8)),
	2776 => std_logic_vector(to_unsigned(173, 8)),
	2777 => std_logic_vector(to_unsigned(173, 8)),
	2778 => std_logic_vector(to_unsigned(163, 8)),
	2779 => std_logic_vector(to_unsigned(169, 8)),
	2780 => std_logic_vector(to_unsigned(169, 8)),
	2781 => std_logic_vector(to_unsigned(164, 8)),
	2782 => std_logic_vector(to_unsigned(171, 8)),
	2783 => std_logic_vector(to_unsigned(175, 8)),
	2784 => std_logic_vector(to_unsigned(167, 8)),
	2785 => std_logic_vector(to_unsigned(167, 8)),
	2786 => std_logic_vector(to_unsigned(171, 8)),
	2787 => std_logic_vector(to_unsigned(162, 8)),
	2788 => std_logic_vector(to_unsigned(163, 8)),
	2789 => std_logic_vector(to_unsigned(169, 8)),
	2790 => std_logic_vector(to_unsigned(166, 8)),
	2791 => std_logic_vector(to_unsigned(163, 8)),
	2792 => std_logic_vector(to_unsigned(166, 8)),
	2793 => std_logic_vector(to_unsigned(171, 8)),
	2794 => std_logic_vector(to_unsigned(169, 8)),
	2795 => std_logic_vector(to_unsigned(166, 8)),
	2796 => std_logic_vector(to_unsigned(170, 8)),
	2797 => std_logic_vector(to_unsigned(172, 8)),
	2798 => std_logic_vector(to_unsigned(172, 8)),
	2799 => std_logic_vector(to_unsigned(162, 8)),
	2800 => std_logic_vector(to_unsigned(176, 8)),
	2801 => std_logic_vector(to_unsigned(168, 8)),
	2802 => std_logic_vector(to_unsigned(172, 8)),
	2803 => std_logic_vector(to_unsigned(176, 8)),
	2804 => std_logic_vector(to_unsigned(170, 8)),
	2805 => std_logic_vector(to_unsigned(169, 8)),
	2806 => std_logic_vector(to_unsigned(173, 8)),
	2807 => std_logic_vector(to_unsigned(176, 8)),
	2808 => std_logic_vector(to_unsigned(166, 8)),
	2809 => std_logic_vector(to_unsigned(166, 8)),
	2810 => std_logic_vector(to_unsigned(167, 8)),
	2811 => std_logic_vector(to_unsigned(171, 8)),
	2812 => std_logic_vector(to_unsigned(164, 8)),
	2813 => std_logic_vector(to_unsigned(173, 8)),
	2814 => std_logic_vector(to_unsigned(171, 8)),
	2815 => std_logic_vector(to_unsigned(163, 8)),
	2816 => std_logic_vector(to_unsigned(165, 8)),
	2817 => std_logic_vector(to_unsigned(163, 8)),
	2818 => std_logic_vector(to_unsigned(169, 8)),
	2819 => std_logic_vector(to_unsigned(162, 8)),
	2820 => std_logic_vector(to_unsigned(163, 8)),
	2821 => std_logic_vector(to_unsigned(163, 8)),
	2822 => std_logic_vector(to_unsigned(174, 8)),
	2823 => std_logic_vector(to_unsigned(171, 8)),
	2824 => std_logic_vector(to_unsigned(168, 8)),
	2825 => std_logic_vector(to_unsigned(176, 8)),
	2826 => std_logic_vector(to_unsigned(169, 8)),
	2827 => std_logic_vector(to_unsigned(162, 8)),
	2828 => std_logic_vector(to_unsigned(166, 8)),
	2829 => std_logic_vector(to_unsigned(171, 8)),
	2830 => std_logic_vector(to_unsigned(172, 8)),
	2831 => std_logic_vector(to_unsigned(168, 8)),
	2832 => std_logic_vector(to_unsigned(173, 8)),
	2833 => std_logic_vector(to_unsigned(175, 8)),
	2834 => std_logic_vector(to_unsigned(162, 8)),
	2835 => std_logic_vector(to_unsigned(173, 8)),
	2836 => std_logic_vector(to_unsigned(171, 8)),
	2837 => std_logic_vector(to_unsigned(175, 8)),
	2838 => std_logic_vector(to_unsigned(170, 8)),
	2839 => std_logic_vector(to_unsigned(162, 8)),
	2840 => std_logic_vector(to_unsigned(174, 8)),
	2841 => std_logic_vector(to_unsigned(165, 8)),
	2842 => std_logic_vector(to_unsigned(176, 8)),
	2843 => std_logic_vector(to_unsigned(163, 8)),
	2844 => std_logic_vector(to_unsigned(165, 8)),
	2845 => std_logic_vector(to_unsigned(164, 8)),
	2846 => std_logic_vector(to_unsigned(163, 8)),
	2847 => std_logic_vector(to_unsigned(174, 8)),
	2848 => std_logic_vector(to_unsigned(172, 8)),
	2849 => std_logic_vector(to_unsigned(168, 8)),
	2850 => std_logic_vector(to_unsigned(176, 8)),
	2851 => std_logic_vector(to_unsigned(163, 8)),
	2852 => std_logic_vector(to_unsigned(172, 8)),
	2853 => std_logic_vector(to_unsigned(162, 8)),
	2854 => std_logic_vector(to_unsigned(174, 8)),
	2855 => std_logic_vector(to_unsigned(163, 8)),
	2856 => std_logic_vector(to_unsigned(166, 8)),
	2857 => std_logic_vector(to_unsigned(175, 8)),
	2858 => std_logic_vector(to_unsigned(176, 8)),
	2859 => std_logic_vector(to_unsigned(175, 8)),
	2860 => std_logic_vector(to_unsigned(175, 8)),
	2861 => std_logic_vector(to_unsigned(165, 8)),
	2862 => std_logic_vector(to_unsigned(163, 8)),
	2863 => std_logic_vector(to_unsigned(176, 8)),
	2864 => std_logic_vector(to_unsigned(165, 8)),
	2865 => std_logic_vector(to_unsigned(166, 8)),
	2866 => std_logic_vector(to_unsigned(172, 8)),
	2867 => std_logic_vector(to_unsigned(171, 8)),
	2868 => std_logic_vector(to_unsigned(164, 8)),
	2869 => std_logic_vector(to_unsigned(170, 8)),
	2870 => std_logic_vector(to_unsigned(162, 8)),
	2871 => std_logic_vector(to_unsigned(176, 8)),
	2872 => std_logic_vector(to_unsigned(166, 8)),
	2873 => std_logic_vector(to_unsigned(173, 8)),
	2874 => std_logic_vector(to_unsigned(175, 8)),
	2875 => std_logic_vector(to_unsigned(169, 8)),
	2876 => std_logic_vector(to_unsigned(168, 8)),
	2877 => std_logic_vector(to_unsigned(166, 8)),
	2878 => std_logic_vector(to_unsigned(165, 8)),
	2879 => std_logic_vector(to_unsigned(166, 8)),
	2880 => std_logic_vector(to_unsigned(162, 8)),
	2881 => std_logic_vector(to_unsigned(162, 8)),
	2882 => std_logic_vector(to_unsigned(176, 8)),
	2883 => std_logic_vector(to_unsigned(162, 8)),
	2884 => std_logic_vector(to_unsigned(162, 8)),
	2885 => std_logic_vector(to_unsigned(171, 8)),
	2886 => std_logic_vector(to_unsigned(175, 8)),
	2887 => std_logic_vector(to_unsigned(162, 8)),
	2888 => std_logic_vector(to_unsigned(167, 8)),
	2889 => std_logic_vector(to_unsigned(175, 8)),
	2890 => std_logic_vector(to_unsigned(172, 8)),
	2891 => std_logic_vector(to_unsigned(173, 8)),
	2892 => std_logic_vector(to_unsigned(167, 8)),
	2893 => std_logic_vector(to_unsigned(172, 8)),
	2894 => std_logic_vector(to_unsigned(168, 8)),
	2895 => std_logic_vector(to_unsigned(162, 8)),
	2896 => std_logic_vector(to_unsigned(166, 8)),
	2897 => std_logic_vector(to_unsigned(169, 8)),
	2898 => std_logic_vector(to_unsigned(176, 8)),
	2899 => std_logic_vector(to_unsigned(164, 8)),
	2900 => std_logic_vector(to_unsigned(176, 8)),
	2901 => std_logic_vector(to_unsigned(173, 8)),
	2902 => std_logic_vector(to_unsigned(167, 8)),
	2903 => std_logic_vector(to_unsigned(171, 8)),
	2904 => std_logic_vector(to_unsigned(175, 8)),
	2905 => std_logic_vector(to_unsigned(172, 8)),
	2906 => std_logic_vector(to_unsigned(173, 8)),
	2907 => std_logic_vector(to_unsigned(165, 8)),
	2908 => std_logic_vector(to_unsigned(169, 8)),
	2909 => std_logic_vector(to_unsigned(176, 8)),
	2910 => std_logic_vector(to_unsigned(174, 8)),
	2911 => std_logic_vector(to_unsigned(165, 8)),
	2912 => std_logic_vector(to_unsigned(169, 8)),
	2913 => std_logic_vector(to_unsigned(164, 8)),
	2914 => std_logic_vector(to_unsigned(164, 8)),
	2915 => std_logic_vector(to_unsigned(171, 8)),
	2916 => std_logic_vector(to_unsigned(169, 8)),
	2917 => std_logic_vector(to_unsigned(164, 8)),
	2918 => std_logic_vector(to_unsigned(176, 8)),
	2919 => std_logic_vector(to_unsigned(170, 8)),
	2920 => std_logic_vector(to_unsigned(175, 8)),
	2921 => std_logic_vector(to_unsigned(175, 8)),
	2922 => std_logic_vector(to_unsigned(172, 8)),
	2923 => std_logic_vector(to_unsigned(174, 8)),
	2924 => std_logic_vector(to_unsigned(169, 8)),
	2925 => std_logic_vector(to_unsigned(170, 8)),
	2926 => std_logic_vector(to_unsigned(166, 8)),
	2927 => std_logic_vector(to_unsigned(173, 8)),
	2928 => std_logic_vector(to_unsigned(170, 8)),
	2929 => std_logic_vector(to_unsigned(174, 8)),
	2930 => std_logic_vector(to_unsigned(172, 8)),
	2931 => std_logic_vector(to_unsigned(162, 8)),
	2932 => std_logic_vector(to_unsigned(169, 8)),
	2933 => std_logic_vector(to_unsigned(168, 8)),
	2934 => std_logic_vector(to_unsigned(163, 8)),
	2935 => std_logic_vector(to_unsigned(168, 8)),
	2936 => std_logic_vector(to_unsigned(165, 8)),
	2937 => std_logic_vector(to_unsigned(173, 8)),
	2938 => std_logic_vector(to_unsigned(176, 8)),
	2939 => std_logic_vector(to_unsigned(163, 8)),
	2940 => std_logic_vector(to_unsigned(164, 8)),
	2941 => std_logic_vector(to_unsigned(175, 8)),
	2942 => std_logic_vector(to_unsigned(172, 8)),
	2943 => std_logic_vector(to_unsigned(168, 8)),
	2944 => std_logic_vector(to_unsigned(172, 8)),
	2945 => std_logic_vector(to_unsigned(167, 8)),
	2946 => std_logic_vector(to_unsigned(165, 8)),
	2947 => std_logic_vector(to_unsigned(165, 8)),
	2948 => std_logic_vector(to_unsigned(169, 8)),
	2949 => std_logic_vector(to_unsigned(167, 8)),
	2950 => std_logic_vector(to_unsigned(173, 8)),
	2951 => std_logic_vector(to_unsigned(168, 8)),
	2952 => std_logic_vector(to_unsigned(168, 8)),
	2953 => std_logic_vector(to_unsigned(162, 8)),
	2954 => std_logic_vector(to_unsigned(165, 8)),
	2955 => std_logic_vector(to_unsigned(171, 8)),
	2956 => std_logic_vector(to_unsigned(174, 8)),
	2957 => std_logic_vector(to_unsigned(166, 8)),
	2958 => std_logic_vector(to_unsigned(172, 8)),
	2959 => std_logic_vector(to_unsigned(169, 8)),
	2960 => std_logic_vector(to_unsigned(169, 8)),
	2961 => std_logic_vector(to_unsigned(166, 8)),
	2962 => std_logic_vector(to_unsigned(167, 8)),
	2963 => std_logic_vector(to_unsigned(176, 8)),
	2964 => std_logic_vector(to_unsigned(169, 8)),
	2965 => std_logic_vector(to_unsigned(169, 8)),
	2966 => std_logic_vector(to_unsigned(171, 8)),
	2967 => std_logic_vector(to_unsigned(164, 8)),
	2968 => std_logic_vector(to_unsigned(167, 8)),
	2969 => std_logic_vector(to_unsigned(167, 8)),
	2970 => std_logic_vector(to_unsigned(162, 8)),
	2971 => std_logic_vector(to_unsigned(170, 8)),
	2972 => std_logic_vector(to_unsigned(162, 8)),
	2973 => std_logic_vector(to_unsigned(162, 8)),
	2974 => std_logic_vector(to_unsigned(175, 8)),
	2975 => std_logic_vector(to_unsigned(163, 8)),
	2976 => std_logic_vector(to_unsigned(171, 8)),
	2977 => std_logic_vector(to_unsigned(175, 8)),
	2978 => std_logic_vector(to_unsigned(163, 8)),
	2979 => std_logic_vector(to_unsigned(169, 8)),
	2980 => std_logic_vector(to_unsigned(175, 8)),
	2981 => std_logic_vector(to_unsigned(164, 8)),
	2982 => std_logic_vector(to_unsigned(168, 8)),
	2983 => std_logic_vector(to_unsigned(162, 8)),
	2984 => std_logic_vector(to_unsigned(166, 8)),
	2985 => std_logic_vector(to_unsigned(173, 8)),
	2986 => std_logic_vector(to_unsigned(176, 8)),
	2987 => std_logic_vector(to_unsigned(175, 8)),
	2988 => std_logic_vector(to_unsigned(165, 8)),
	2989 => std_logic_vector(to_unsigned(171, 8)),
	2990 => std_logic_vector(to_unsigned(173, 8)),
	2991 => std_logic_vector(to_unsigned(176, 8)),
	2992 => std_logic_vector(to_unsigned(163, 8)),
	2993 => std_logic_vector(to_unsigned(175, 8)),
	2994 => std_logic_vector(to_unsigned(174, 8)),
	2995 => std_logic_vector(to_unsigned(172, 8)),
	2996 => std_logic_vector(to_unsigned(166, 8)),
	2997 => std_logic_vector(to_unsigned(171, 8)),
	2998 => std_logic_vector(to_unsigned(170, 8)),
	2999 => std_logic_vector(to_unsigned(165, 8)),
	3000 => std_logic_vector(to_unsigned(164, 8)),
	3001 => std_logic_vector(to_unsigned(173, 8)),
	3002 => std_logic_vector(to_unsigned(170, 8)),
	3003 => std_logic_vector(to_unsigned(164, 8)),
	3004 => std_logic_vector(to_unsigned(165, 8)),
	3005 => std_logic_vector(to_unsigned(174, 8)),
	3006 => std_logic_vector(to_unsigned(164, 8)),
	3007 => std_logic_vector(to_unsigned(162, 8)),
	3008 => std_logic_vector(to_unsigned(166, 8)),
	3009 => std_logic_vector(to_unsigned(165, 8)),
	3010 => std_logic_vector(to_unsigned(168, 8)),
	3011 => std_logic_vector(to_unsigned(166, 8)),
	3012 => std_logic_vector(to_unsigned(164, 8)),
	3013 => std_logic_vector(to_unsigned(164, 8)),
	3014 => std_logic_vector(to_unsigned(173, 8)),
	3015 => std_logic_vector(to_unsigned(168, 8)),
	3016 => std_logic_vector(to_unsigned(163, 8)),
	3017 => std_logic_vector(to_unsigned(173, 8)),
	3018 => std_logic_vector(to_unsigned(164, 8)),
	3019 => std_logic_vector(to_unsigned(164, 8)),
	3020 => std_logic_vector(to_unsigned(162, 8)),
	3021 => std_logic_vector(to_unsigned(175, 8)),
	3022 => std_logic_vector(to_unsigned(163, 8)),
	3023 => std_logic_vector(to_unsigned(176, 8)),
	3024 => std_logic_vector(to_unsigned(172, 8)),
	3025 => std_logic_vector(to_unsigned(168, 8)),
	3026 => std_logic_vector(to_unsigned(166, 8)),
	3027 => std_logic_vector(to_unsigned(166, 8)),
	3028 => std_logic_vector(to_unsigned(175, 8)),
	3029 => std_logic_vector(to_unsigned(166, 8)),
	3030 => std_logic_vector(to_unsigned(174, 8)),
	3031 => std_logic_vector(to_unsigned(175, 8)),
	3032 => std_logic_vector(to_unsigned(170, 8)),
	3033 => std_logic_vector(to_unsigned(167, 8)),
	3034 => std_logic_vector(to_unsigned(163, 8)),
	3035 => std_logic_vector(to_unsigned(174, 8)),
	3036 => std_logic_vector(to_unsigned(164, 8)),
	3037 => std_logic_vector(to_unsigned(167, 8)),
	3038 => std_logic_vector(to_unsigned(173, 8)),
	3039 => std_logic_vector(to_unsigned(169, 8)),
	3040 => std_logic_vector(to_unsigned(171, 8)),
	3041 => std_logic_vector(to_unsigned(175, 8)),
	3042 => std_logic_vector(to_unsigned(171, 8)),
	3043 => std_logic_vector(to_unsigned(170, 8)),
	3044 => std_logic_vector(to_unsigned(170, 8)),
	3045 => std_logic_vector(to_unsigned(174, 8)),
	3046 => std_logic_vector(to_unsigned(165, 8)),
	3047 => std_logic_vector(to_unsigned(164, 8)),
	3048 => std_logic_vector(to_unsigned(167, 8)),
	3049 => std_logic_vector(to_unsigned(167, 8)),
	3050 => std_logic_vector(to_unsigned(174, 8)),
	3051 => std_logic_vector(to_unsigned(167, 8)),
	3052 => std_logic_vector(to_unsigned(165, 8)),
	3053 => std_logic_vector(to_unsigned(172, 8)),
	3054 => std_logic_vector(to_unsigned(163, 8)),
	3055 => std_logic_vector(to_unsigned(174, 8)),
	3056 => std_logic_vector(to_unsigned(162, 8)),
	3057 => std_logic_vector(to_unsigned(176, 8)),
	3058 => std_logic_vector(to_unsigned(170, 8)),
	3059 => std_logic_vector(to_unsigned(168, 8)),
	3060 => std_logic_vector(to_unsigned(172, 8)),
	3061 => std_logic_vector(to_unsigned(171, 8)),
	3062 => std_logic_vector(to_unsigned(169, 8)),
	3063 => std_logic_vector(to_unsigned(176, 8)),
	3064 => std_logic_vector(to_unsigned(176, 8)),
	3065 => std_logic_vector(to_unsigned(171, 8)),
	3066 => std_logic_vector(to_unsigned(170, 8)),
	3067 => std_logic_vector(to_unsigned(169, 8)),
	3068 => std_logic_vector(to_unsigned(170, 8)),
	3069 => std_logic_vector(to_unsigned(164, 8)),
	3070 => std_logic_vector(to_unsigned(162, 8)),
	3071 => std_logic_vector(to_unsigned(174, 8)),
	3072 => std_logic_vector(to_unsigned(165, 8)),
	3073 => std_logic_vector(to_unsigned(169, 8)),
	3074 => std_logic_vector(to_unsigned(176, 8)),
	3075 => std_logic_vector(to_unsigned(163, 8)),
	3076 => std_logic_vector(to_unsigned(173, 8)),
	3077 => std_logic_vector(to_unsigned(171, 8)),
	3078 => std_logic_vector(to_unsigned(173, 8)),
	3079 => std_logic_vector(to_unsigned(166, 8)),
	3080 => std_logic_vector(to_unsigned(176, 8)),
	3081 => std_logic_vector(to_unsigned(163, 8)),
	3082 => std_logic_vector(to_unsigned(175, 8)),
	3083 => std_logic_vector(to_unsigned(169, 8)),
	3084 => std_logic_vector(to_unsigned(173, 8)),
	3085 => std_logic_vector(to_unsigned(169, 8)),
	3086 => std_logic_vector(to_unsigned(172, 8)),
	3087 => std_logic_vector(to_unsigned(163, 8)),
	3088 => std_logic_vector(to_unsigned(176, 8)),
	3089 => std_logic_vector(to_unsigned(172, 8)),
	3090 => std_logic_vector(to_unsigned(168, 8)),
	3091 => std_logic_vector(to_unsigned(165, 8)),
	3092 => std_logic_vector(to_unsigned(168, 8)),
	3093 => std_logic_vector(to_unsigned(165, 8)),
	3094 => std_logic_vector(to_unsigned(165, 8)),
	3095 => std_logic_vector(to_unsigned(165, 8)),
	3096 => std_logic_vector(to_unsigned(171, 8)),
	3097 => std_logic_vector(to_unsigned(176, 8)),
	3098 => std_logic_vector(to_unsigned(170, 8)),
	3099 => std_logic_vector(to_unsigned(168, 8)),
	3100 => std_logic_vector(to_unsigned(164, 8)),
	3101 => std_logic_vector(to_unsigned(162, 8)),
	3102 => std_logic_vector(to_unsigned(175, 8)),
	3103 => std_logic_vector(to_unsigned(171, 8)),
	3104 => std_logic_vector(to_unsigned(166, 8)),
	3105 => std_logic_vector(to_unsigned(162, 8)),
	3106 => std_logic_vector(to_unsigned(169, 8)),
	3107 => std_logic_vector(to_unsigned(163, 8)),
	3108 => std_logic_vector(to_unsigned(172, 8)),
	3109 => std_logic_vector(to_unsigned(166, 8)),
	3110 => std_logic_vector(to_unsigned(176, 8)),
	3111 => std_logic_vector(to_unsigned(168, 8)),
	3112 => std_logic_vector(to_unsigned(167, 8)),
	3113 => std_logic_vector(to_unsigned(169, 8)),
	3114 => std_logic_vector(to_unsigned(166, 8)),
	3115 => std_logic_vector(to_unsigned(174, 8)),
	3116 => std_logic_vector(to_unsigned(175, 8)),
	3117 => std_logic_vector(to_unsigned(170, 8)),
	3118 => std_logic_vector(to_unsigned(172, 8)),
	3119 => std_logic_vector(to_unsigned(173, 8)),
	3120 => std_logic_vector(to_unsigned(174, 8)),
	3121 => std_logic_vector(to_unsigned(170, 8)),
	3122 => std_logic_vector(to_unsigned(167, 8)),
	3123 => std_logic_vector(to_unsigned(172, 8)),
	3124 => std_logic_vector(to_unsigned(172, 8)),
	3125 => std_logic_vector(to_unsigned(171, 8)),
	3126 => std_logic_vector(to_unsigned(173, 8)),
	3127 => std_logic_vector(to_unsigned(162, 8)),
	3128 => std_logic_vector(to_unsigned(166, 8)),
	3129 => std_logic_vector(to_unsigned(165, 8)),
	3130 => std_logic_vector(to_unsigned(176, 8)),
	3131 => std_logic_vector(to_unsigned(164, 8)),
	3132 => std_logic_vector(to_unsigned(168, 8)),
	3133 => std_logic_vector(to_unsigned(165, 8)),
	3134 => std_logic_vector(to_unsigned(164, 8)),
	3135 => std_logic_vector(to_unsigned(165, 8)),
	3136 => std_logic_vector(to_unsigned(163, 8)),
	3137 => std_logic_vector(to_unsigned(162, 8)),
	3138 => std_logic_vector(to_unsigned(163, 8)),
	3139 => std_logic_vector(to_unsigned(166, 8)),
	3140 => std_logic_vector(to_unsigned(162, 8)),
	3141 => std_logic_vector(to_unsigned(171, 8)),
	3142 => std_logic_vector(to_unsigned(162, 8)),
	3143 => std_logic_vector(to_unsigned(174, 8)),
	3144 => std_logic_vector(to_unsigned(169, 8)),
	3145 => std_logic_vector(to_unsigned(162, 8)),
	3146 => std_logic_vector(to_unsigned(171, 8)),
	3147 => std_logic_vector(to_unsigned(176, 8)),
	3148 => std_logic_vector(to_unsigned(174, 8)),
	3149 => std_logic_vector(to_unsigned(166, 8)),
	3150 => std_logic_vector(to_unsigned(166, 8)),
	3151 => std_logic_vector(to_unsigned(166, 8)),
	3152 => std_logic_vector(to_unsigned(162, 8)),
	3153 => std_logic_vector(to_unsigned(165, 8)),
	3154 => std_logic_vector(to_unsigned(164, 8)),
	3155 => std_logic_vector(to_unsigned(167, 8)),
	3156 => std_logic_vector(to_unsigned(162, 8)),
	3157 => std_logic_vector(to_unsigned(170, 8)),
	3158 => std_logic_vector(to_unsigned(170, 8)),
	3159 => std_logic_vector(to_unsigned(166, 8)),
	3160 => std_logic_vector(to_unsigned(167, 8)),
	3161 => std_logic_vector(to_unsigned(176, 8)),
	3162 => std_logic_vector(to_unsigned(175, 8)),
	3163 => std_logic_vector(to_unsigned(175, 8)),
	3164 => std_logic_vector(to_unsigned(166, 8)),
	3165 => std_logic_vector(to_unsigned(163, 8)),
	3166 => std_logic_vector(to_unsigned(169, 8)),
	3167 => std_logic_vector(to_unsigned(162, 8)),
	3168 => std_logic_vector(to_unsigned(174, 8)),
	3169 => std_logic_vector(to_unsigned(167, 8)),
	3170 => std_logic_vector(to_unsigned(176, 8)),
	3171 => std_logic_vector(to_unsigned(165, 8)),
	3172 => std_logic_vector(to_unsigned(169, 8)),
	3173 => std_logic_vector(to_unsigned(165, 8)),
	3174 => std_logic_vector(to_unsigned(170, 8)),
	3175 => std_logic_vector(to_unsigned(170, 8)),
	3176 => std_logic_vector(to_unsigned(173, 8)),
	3177 => std_logic_vector(to_unsigned(170, 8)),
	3178 => std_logic_vector(to_unsigned(174, 8)),
	3179 => std_logic_vector(to_unsigned(167, 8)),
	3180 => std_logic_vector(to_unsigned(164, 8)),
	3181 => std_logic_vector(to_unsigned(176, 8)),
	3182 => std_logic_vector(to_unsigned(168, 8)),
	3183 => std_logic_vector(to_unsigned(167, 8)),
	3184 => std_logic_vector(to_unsigned(169, 8)),
	3185 => std_logic_vector(to_unsigned(167, 8)),
	3186 => std_logic_vector(to_unsigned(163, 8)),
	3187 => std_logic_vector(to_unsigned(167, 8)),
	3188 => std_logic_vector(to_unsigned(162, 8)),
	3189 => std_logic_vector(to_unsigned(168, 8)),
	3190 => std_logic_vector(to_unsigned(172, 8)),
	3191 => std_logic_vector(to_unsigned(176, 8)),
	3192 => std_logic_vector(to_unsigned(168, 8)),
	3193 => std_logic_vector(to_unsigned(163, 8)),
	3194 => std_logic_vector(to_unsigned(170, 8)),
	3195 => std_logic_vector(to_unsigned(170, 8)),
	3196 => std_logic_vector(to_unsigned(168, 8)),
	3197 => std_logic_vector(to_unsigned(174, 8)),
	3198 => std_logic_vector(to_unsigned(176, 8)),
	3199 => std_logic_vector(to_unsigned(162, 8)),
	3200 => std_logic_vector(to_unsigned(166, 8)),
	3201 => std_logic_vector(to_unsigned(171, 8)),
	3202 => std_logic_vector(to_unsigned(164, 8)),
	3203 => std_logic_vector(to_unsigned(163, 8)),
	3204 => std_logic_vector(to_unsigned(163, 8)),
	3205 => std_logic_vector(to_unsigned(170, 8)),
	3206 => std_logic_vector(to_unsigned(173, 8)),
	3207 => std_logic_vector(to_unsigned(166, 8)),
	3208 => std_logic_vector(to_unsigned(173, 8)),
	3209 => std_logic_vector(to_unsigned(175, 8)),
	3210 => std_logic_vector(to_unsigned(164, 8)),
	3211 => std_logic_vector(to_unsigned(172, 8)),
	3212 => std_logic_vector(to_unsigned(166, 8)),
	3213 => std_logic_vector(to_unsigned(173, 8)),
	3214 => std_logic_vector(to_unsigned(169, 8)),
	3215 => std_logic_vector(to_unsigned(169, 8)),
	3216 => std_logic_vector(to_unsigned(171, 8)),
	3217 => std_logic_vector(to_unsigned(174, 8)),
	3218 => std_logic_vector(to_unsigned(170, 8)),
	3219 => std_logic_vector(to_unsigned(173, 8)),
	3220 => std_logic_vector(to_unsigned(175, 8)),
	3221 => std_logic_vector(to_unsigned(175, 8)),
	3222 => std_logic_vector(to_unsigned(168, 8)),
	3223 => std_logic_vector(to_unsigned(170, 8)),
	3224 => std_logic_vector(to_unsigned(170, 8)),
	3225 => std_logic_vector(to_unsigned(169, 8)),
	3226 => std_logic_vector(to_unsigned(170, 8)),
	3227 => std_logic_vector(to_unsigned(175, 8)),
	3228 => std_logic_vector(to_unsigned(167, 8)),
	3229 => std_logic_vector(to_unsigned(165, 8)),
	3230 => std_logic_vector(to_unsigned(165, 8)),
	3231 => std_logic_vector(to_unsigned(173, 8)),
	3232 => std_logic_vector(to_unsigned(172, 8)),
	3233 => std_logic_vector(to_unsigned(168, 8)),
	3234 => std_logic_vector(to_unsigned(172, 8)),
	3235 => std_logic_vector(to_unsigned(167, 8)),
	3236 => std_logic_vector(to_unsigned(171, 8)),
	3237 => std_logic_vector(to_unsigned(172, 8)),
	3238 => std_logic_vector(to_unsigned(169, 8)),
	3239 => std_logic_vector(to_unsigned(168, 8)),
	3240 => std_logic_vector(to_unsigned(167, 8)),
	3241 => std_logic_vector(to_unsigned(176, 8)),
	3242 => std_logic_vector(to_unsigned(168, 8)),
	3243 => std_logic_vector(to_unsigned(172, 8)),
	3244 => std_logic_vector(to_unsigned(172, 8)),
	3245 => std_logic_vector(to_unsigned(168, 8)),
	3246 => std_logic_vector(to_unsigned(176, 8)),
	3247 => std_logic_vector(to_unsigned(173, 8)),
	3248 => std_logic_vector(to_unsigned(163, 8)),
	3249 => std_logic_vector(to_unsigned(169, 8)),
	3250 => std_logic_vector(to_unsigned(174, 8)),
	3251 => std_logic_vector(to_unsigned(171, 8)),
	3252 => std_logic_vector(to_unsigned(168, 8)),
	3253 => std_logic_vector(to_unsigned(176, 8)),
	3254 => std_logic_vector(to_unsigned(170, 8)),
	3255 => std_logic_vector(to_unsigned(172, 8)),
	3256 => std_logic_vector(to_unsigned(163, 8)),
	3257 => std_logic_vector(to_unsigned(171, 8)),
	3258 => std_logic_vector(to_unsigned(170, 8)),
	3259 => std_logic_vector(to_unsigned(165, 8)),
	3260 => std_logic_vector(to_unsigned(174, 8)),
	3261 => std_logic_vector(to_unsigned(172, 8)),
	3262 => std_logic_vector(to_unsigned(172, 8)),
	3263 => std_logic_vector(to_unsigned(173, 8)),
	3264 => std_logic_vector(to_unsigned(164, 8)),
	3265 => std_logic_vector(to_unsigned(173, 8)),
	3266 => std_logic_vector(to_unsigned(175, 8)),
	3267 => std_logic_vector(to_unsigned(163, 8)),
	3268 => std_logic_vector(to_unsigned(165, 8)),
	3269 => std_logic_vector(to_unsigned(167, 8)),
	3270 => std_logic_vector(to_unsigned(163, 8)),
	3271 => std_logic_vector(to_unsigned(162, 8)),
	3272 => std_logic_vector(to_unsigned(174, 8)),
	3273 => std_logic_vector(to_unsigned(163, 8)),
	3274 => std_logic_vector(to_unsigned(172, 8)),
	3275 => std_logic_vector(to_unsigned(165, 8)),
	3276 => std_logic_vector(to_unsigned(162, 8)),
	3277 => std_logic_vector(to_unsigned(169, 8)),
	3278 => std_logic_vector(to_unsigned(167, 8)),
	3279 => std_logic_vector(to_unsigned(167, 8)),
	3280 => std_logic_vector(to_unsigned(172, 8)),
	3281 => std_logic_vector(to_unsigned(173, 8)),
	3282 => std_logic_vector(to_unsigned(174, 8)),
	3283 => std_logic_vector(to_unsigned(166, 8)),
	3284 => std_logic_vector(to_unsigned(167, 8)),
	3285 => std_logic_vector(to_unsigned(171, 8)),
	3286 => std_logic_vector(to_unsigned(169, 8)),
	3287 => std_logic_vector(to_unsigned(164, 8)),
	3288 => std_logic_vector(to_unsigned(170, 8)),
	3289 => std_logic_vector(to_unsigned(174, 8)),
	3290 => std_logic_vector(to_unsigned(175, 8)),
	3291 => std_logic_vector(to_unsigned(170, 8)),
	3292 => std_logic_vector(to_unsigned(172, 8)),
	3293 => std_logic_vector(to_unsigned(174, 8)),
	3294 => std_logic_vector(to_unsigned(167, 8)),
	3295 => std_logic_vector(to_unsigned(168, 8)),
	3296 => std_logic_vector(to_unsigned(171, 8)),
	3297 => std_logic_vector(to_unsigned(174, 8)),
	3298 => std_logic_vector(to_unsigned(174, 8)),
	3299 => std_logic_vector(to_unsigned(164, 8)),
	3300 => std_logic_vector(to_unsigned(164, 8)),
	3301 => std_logic_vector(to_unsigned(173, 8)),
	3302 => std_logic_vector(to_unsigned(175, 8)),
	3303 => std_logic_vector(to_unsigned(169, 8)),
	3304 => std_logic_vector(to_unsigned(176, 8)),
	3305 => std_logic_vector(to_unsigned(168, 8)),
	3306 => std_logic_vector(to_unsigned(165, 8)),
	3307 => std_logic_vector(to_unsigned(167, 8)),
	3308 => std_logic_vector(to_unsigned(175, 8)),
	3309 => std_logic_vector(to_unsigned(169, 8)),
	3310 => std_logic_vector(to_unsigned(174, 8)),
	3311 => std_logic_vector(to_unsigned(171, 8)),
	3312 => std_logic_vector(to_unsigned(171, 8)),
	3313 => std_logic_vector(to_unsigned(166, 8)),
	3314 => std_logic_vector(to_unsigned(167, 8)),
	3315 => std_logic_vector(to_unsigned(164, 8)),
	3316 => std_logic_vector(to_unsigned(163, 8)),
	3317 => std_logic_vector(to_unsigned(174, 8)),
	3318 => std_logic_vector(to_unsigned(165, 8)),
	3319 => std_logic_vector(to_unsigned(170, 8)),
	3320 => std_logic_vector(to_unsigned(168, 8)),
	3321 => std_logic_vector(to_unsigned(169, 8)),
	3322 => std_logic_vector(to_unsigned(174, 8)),
	3323 => std_logic_vector(to_unsigned(168, 8)),
	3324 => std_logic_vector(to_unsigned(167, 8)),
	3325 => std_logic_vector(to_unsigned(168, 8)),
	3326 => std_logic_vector(to_unsigned(165, 8)),
	3327 => std_logic_vector(to_unsigned(171, 8)),
	3328 => std_logic_vector(to_unsigned(170, 8)),
	3329 => std_logic_vector(to_unsigned(167, 8)),
	3330 => std_logic_vector(to_unsigned(162, 8)),
	3331 => std_logic_vector(to_unsigned(166, 8)),
	3332 => std_logic_vector(to_unsigned(176, 8)),
	3333 => std_logic_vector(to_unsigned(169, 8)),
	3334 => std_logic_vector(to_unsigned(173, 8)),
	3335 => std_logic_vector(to_unsigned(172, 8)),
	3336 => std_logic_vector(to_unsigned(162, 8)),
	3337 => std_logic_vector(to_unsigned(165, 8)),
	3338 => std_logic_vector(to_unsigned(165, 8)),
	3339 => std_logic_vector(to_unsigned(172, 8)),
	3340 => std_logic_vector(to_unsigned(165, 8)),
	3341 => std_logic_vector(to_unsigned(170, 8)),
	3342 => std_logic_vector(to_unsigned(175, 8)),
	3343 => std_logic_vector(to_unsigned(174, 8)),
	3344 => std_logic_vector(to_unsigned(167, 8)),
	3345 => std_logic_vector(to_unsigned(163, 8)),
	3346 => std_logic_vector(to_unsigned(173, 8)),
	3347 => std_logic_vector(to_unsigned(162, 8)),
	3348 => std_logic_vector(to_unsigned(163, 8)),
	3349 => std_logic_vector(to_unsigned(164, 8)),
	3350 => std_logic_vector(to_unsigned(169, 8)),
	3351 => std_logic_vector(to_unsigned(171, 8)),
	3352 => std_logic_vector(to_unsigned(163, 8)),
	3353 => std_logic_vector(to_unsigned(176, 8)),
	3354 => std_logic_vector(to_unsigned(176, 8)),
	3355 => std_logic_vector(to_unsigned(162, 8)),
	3356 => std_logic_vector(to_unsigned(170, 8)),
	3357 => std_logic_vector(to_unsigned(170, 8)),
	3358 => std_logic_vector(to_unsigned(166, 8)),
	3359 => std_logic_vector(to_unsigned(167, 8)),
	3360 => std_logic_vector(to_unsigned(172, 8)),
	3361 => std_logic_vector(to_unsigned(168, 8)),
	3362 => std_logic_vector(to_unsigned(165, 8)),
	3363 => std_logic_vector(to_unsigned(164, 8)),
	3364 => std_logic_vector(to_unsigned(171, 8)),
	3365 => std_logic_vector(to_unsigned(165, 8)),
	3366 => std_logic_vector(to_unsigned(169, 8)),
	3367 => std_logic_vector(to_unsigned(174, 8)),
	3368 => std_logic_vector(to_unsigned(169, 8)),
	3369 => std_logic_vector(to_unsigned(165, 8)),
	3370 => std_logic_vector(to_unsigned(165, 8)),
	3371 => std_logic_vector(to_unsigned(169, 8)),
	3372 => std_logic_vector(to_unsigned(168, 8)),
	3373 => std_logic_vector(to_unsigned(165, 8)),
	3374 => std_logic_vector(to_unsigned(167, 8)),
	3375 => std_logic_vector(to_unsigned(171, 8)),
	3376 => std_logic_vector(to_unsigned(171, 8)),
	3377 => std_logic_vector(to_unsigned(173, 8)),
	3378 => std_logic_vector(to_unsigned(176, 8)),
	3379 => std_logic_vector(to_unsigned(167, 8)),
	3380 => std_logic_vector(to_unsigned(162, 8)),
	3381 => std_logic_vector(to_unsigned(175, 8)),
	3382 => std_logic_vector(to_unsigned(174, 8)),
	3383 => std_logic_vector(to_unsigned(172, 8)),
	3384 => std_logic_vector(to_unsigned(164, 8)),
	3385 => std_logic_vector(to_unsigned(166, 8)),
	3386 => std_logic_vector(to_unsigned(171, 8)),
	3387 => std_logic_vector(to_unsigned(165, 8)),
	3388 => std_logic_vector(to_unsigned(165, 8)),
	3389 => std_logic_vector(to_unsigned(162, 8)),
	3390 => std_logic_vector(to_unsigned(163, 8)),
	3391 => std_logic_vector(to_unsigned(169, 8)),
	3392 => std_logic_vector(to_unsigned(166, 8)),
	3393 => std_logic_vector(to_unsigned(166, 8)),
	3394 => std_logic_vector(to_unsigned(166, 8)),
	3395 => std_logic_vector(to_unsigned(163, 8)),
	3396 => std_logic_vector(to_unsigned(171, 8)),
	3397 => std_logic_vector(to_unsigned(175, 8)),
	3398 => std_logic_vector(to_unsigned(175, 8)),
	3399 => std_logic_vector(to_unsigned(173, 8)),
	3400 => std_logic_vector(to_unsigned(163, 8)),
	3401 => std_logic_vector(to_unsigned(163, 8)),
	3402 => std_logic_vector(to_unsigned(167, 8)),
	3403 => std_logic_vector(to_unsigned(173, 8)),
	3404 => std_logic_vector(to_unsigned(171, 8)),
	3405 => std_logic_vector(to_unsigned(166, 8)),
	3406 => std_logic_vector(to_unsigned(172, 8)),
	3407 => std_logic_vector(to_unsigned(176, 8)),
	3408 => std_logic_vector(to_unsigned(166, 8)),
	3409 => std_logic_vector(to_unsigned(173, 8)),
	3410 => std_logic_vector(to_unsigned(170, 8)),
	3411 => std_logic_vector(to_unsigned(175, 8)),
	3412 => std_logic_vector(to_unsigned(164, 8)),
	3413 => std_logic_vector(to_unsigned(164, 8)),
	3414 => std_logic_vector(to_unsigned(171, 8)),
	3415 => std_logic_vector(to_unsigned(169, 8)),
	3416 => std_logic_vector(to_unsigned(169, 8)),
	3417 => std_logic_vector(to_unsigned(166, 8)),
	3418 => std_logic_vector(to_unsigned(176, 8)),
	3419 => std_logic_vector(to_unsigned(175, 8)),
	3420 => std_logic_vector(to_unsigned(167, 8)),
	3421 => std_logic_vector(to_unsigned(173, 8)),
	3422 => std_logic_vector(to_unsigned(173, 8)),
	3423 => std_logic_vector(to_unsigned(164, 8)),
	3424 => std_logic_vector(to_unsigned(170, 8)),
	3425 => std_logic_vector(to_unsigned(176, 8)),
	3426 => std_logic_vector(to_unsigned(174, 8)),
	3427 => std_logic_vector(to_unsigned(173, 8)),
	3428 => std_logic_vector(to_unsigned(173, 8)),
	3429 => std_logic_vector(to_unsigned(168, 8)),
	3430 => std_logic_vector(to_unsigned(174, 8)),
	3431 => std_logic_vector(to_unsigned(174, 8)),
	3432 => std_logic_vector(to_unsigned(172, 8)),
	3433 => std_logic_vector(to_unsigned(172, 8)),
	3434 => std_logic_vector(to_unsigned(165, 8)),
	3435 => std_logic_vector(to_unsigned(168, 8)),
	3436 => std_logic_vector(to_unsigned(175, 8)),
	3437 => std_logic_vector(to_unsigned(163, 8)),
	3438 => std_logic_vector(to_unsigned(171, 8)),
	3439 => std_logic_vector(to_unsigned(174, 8)),
	3440 => std_logic_vector(to_unsigned(173, 8)),
	3441 => std_logic_vector(to_unsigned(166, 8)),
	3442 => std_logic_vector(to_unsigned(169, 8)),
	3443 => std_logic_vector(to_unsigned(173, 8)),
	3444 => std_logic_vector(to_unsigned(166, 8)),
	3445 => std_logic_vector(to_unsigned(168, 8)),
	3446 => std_logic_vector(to_unsigned(175, 8)),
	3447 => std_logic_vector(to_unsigned(164, 8)),
	3448 => std_logic_vector(to_unsigned(167, 8)),
	3449 => std_logic_vector(to_unsigned(176, 8)),
	3450 => std_logic_vector(to_unsigned(165, 8)),
	3451 => std_logic_vector(to_unsigned(168, 8)),
	3452 => std_logic_vector(to_unsigned(171, 8)),
	3453 => std_logic_vector(to_unsigned(172, 8)),
	3454 => std_logic_vector(to_unsigned(164, 8)),
	3455 => std_logic_vector(to_unsigned(174, 8)),
	3456 => std_logic_vector(to_unsigned(166, 8)),
	3457 => std_logic_vector(to_unsigned(162, 8)),
	3458 => std_logic_vector(to_unsigned(173, 8)),
	3459 => std_logic_vector(to_unsigned(170, 8)),
	3460 => std_logic_vector(to_unsigned(162, 8)),
	3461 => std_logic_vector(to_unsigned(173, 8)),
	3462 => std_logic_vector(to_unsigned(163, 8)),
	3463 => std_logic_vector(to_unsigned(170, 8)),
	3464 => std_logic_vector(to_unsigned(174, 8)),
	3465 => std_logic_vector(to_unsigned(166, 8)),
	3466 => std_logic_vector(to_unsigned(175, 8)),
	3467 => std_logic_vector(to_unsigned(172, 8)),
	3468 => std_logic_vector(to_unsigned(164, 8)),
	3469 => std_logic_vector(to_unsigned(165, 8)),
	3470 => std_logic_vector(to_unsigned(168, 8)),
	3471 => std_logic_vector(to_unsigned(172, 8)),
	3472 => std_logic_vector(to_unsigned(165, 8)),
	3473 => std_logic_vector(to_unsigned(162, 8)),
	3474 => std_logic_vector(to_unsigned(162, 8)),
	3475 => std_logic_vector(to_unsigned(163, 8)),
	3476 => std_logic_vector(to_unsigned(175, 8)),
	3477 => std_logic_vector(to_unsigned(165, 8)),
	3478 => std_logic_vector(to_unsigned(173, 8)),
	3479 => std_logic_vector(to_unsigned(172, 8)),
	3480 => std_logic_vector(to_unsigned(163, 8)),
	3481 => std_logic_vector(to_unsigned(164, 8)),
	3482 => std_logic_vector(to_unsigned(176, 8)),
	3483 => std_logic_vector(to_unsigned(176, 8)),
	3484 => std_logic_vector(to_unsigned(167, 8)),
	3485 => std_logic_vector(to_unsigned(170, 8)),
	3486 => std_logic_vector(to_unsigned(165, 8)),
	3487 => std_logic_vector(to_unsigned(169, 8)),
	3488 => std_logic_vector(to_unsigned(169, 8)),
	3489 => std_logic_vector(to_unsigned(175, 8)),
	3490 => std_logic_vector(to_unsigned(176, 8)),
	3491 => std_logic_vector(to_unsigned(167, 8)),
	3492 => std_logic_vector(to_unsigned(173, 8)),
	3493 => std_logic_vector(to_unsigned(165, 8)),
	3494 => std_logic_vector(to_unsigned(171, 8)),
	3495 => std_logic_vector(to_unsigned(166, 8)),
	3496 => std_logic_vector(to_unsigned(175, 8)),
	3497 => std_logic_vector(to_unsigned(176, 8)),
	3498 => std_logic_vector(to_unsigned(167, 8)),
	3499 => std_logic_vector(to_unsigned(165, 8)),
	3500 => std_logic_vector(to_unsigned(162, 8)),
	3501 => std_logic_vector(to_unsigned(165, 8)),
	3502 => std_logic_vector(to_unsigned(163, 8)),
	3503 => std_logic_vector(to_unsigned(166, 8)),
	3504 => std_logic_vector(to_unsigned(174, 8)),
	3505 => std_logic_vector(to_unsigned(163, 8)),
	3506 => std_logic_vector(to_unsigned(168, 8)),
	3507 => std_logic_vector(to_unsigned(168, 8)),
	3508 => std_logic_vector(to_unsigned(174, 8)),
	3509 => std_logic_vector(to_unsigned(174, 8)),
	3510 => std_logic_vector(to_unsigned(174, 8)),
	3511 => std_logic_vector(to_unsigned(163, 8)),
	3512 => std_logic_vector(to_unsigned(168, 8)),
	3513 => std_logic_vector(to_unsigned(172, 8)),
	3514 => std_logic_vector(to_unsigned(166, 8)),
	3515 => std_logic_vector(to_unsigned(164, 8)),
	3516 => std_logic_vector(to_unsigned(169, 8)),
	3517 => std_logic_vector(to_unsigned(170, 8)),
	3518 => std_logic_vector(to_unsigned(176, 8)),
	3519 => std_logic_vector(to_unsigned(172, 8)),
	3520 => std_logic_vector(to_unsigned(162, 8)),
	3521 => std_logic_vector(to_unsigned(170, 8)),
	3522 => std_logic_vector(to_unsigned(168, 8)),
	3523 => std_logic_vector(to_unsigned(171, 8)),
	3524 => std_logic_vector(to_unsigned(168, 8)),
	3525 => std_logic_vector(to_unsigned(166, 8)),
	3526 => std_logic_vector(to_unsigned(174, 8)),
	3527 => std_logic_vector(to_unsigned(171, 8)),
	3528 => std_logic_vector(to_unsigned(174, 8)),
	3529 => std_logic_vector(to_unsigned(169, 8)),
	3530 => std_logic_vector(to_unsigned(175, 8)),
	3531 => std_logic_vector(to_unsigned(162, 8)),
	3532 => std_logic_vector(to_unsigned(167, 8)),
	3533 => std_logic_vector(to_unsigned(170, 8)),
	3534 => std_logic_vector(to_unsigned(168, 8)),
	3535 => std_logic_vector(to_unsigned(164, 8)),
	3536 => std_logic_vector(to_unsigned(170, 8)),
	3537 => std_logic_vector(to_unsigned(163, 8)),
	3538 => std_logic_vector(to_unsigned(165, 8)),
	3539 => std_logic_vector(to_unsigned(170, 8)),
	3540 => std_logic_vector(to_unsigned(162, 8)),
	3541 => std_logic_vector(to_unsigned(170, 8)),
	3542 => std_logic_vector(to_unsigned(168, 8)),
	3543 => std_logic_vector(to_unsigned(176, 8)),
	3544 => std_logic_vector(to_unsigned(169, 8)),
	3545 => std_logic_vector(to_unsigned(170, 8)),
	3546 => std_logic_vector(to_unsigned(173, 8)),
	3547 => std_logic_vector(to_unsigned(164, 8)),
	3548 => std_logic_vector(to_unsigned(165, 8)),
	3549 => std_logic_vector(to_unsigned(172, 8)),
	3550 => std_logic_vector(to_unsigned(172, 8)),
	3551 => std_logic_vector(to_unsigned(166, 8)),
	3552 => std_logic_vector(to_unsigned(170, 8)),
	3553 => std_logic_vector(to_unsigned(170, 8)),
	3554 => std_logic_vector(to_unsigned(164, 8)),
	3555 => std_logic_vector(to_unsigned(163, 8)),
	3556 => std_logic_vector(to_unsigned(171, 8)),
	3557 => std_logic_vector(to_unsigned(170, 8)),
	3558 => std_logic_vector(to_unsigned(165, 8)),
	3559 => std_logic_vector(to_unsigned(175, 8)),
	3560 => std_logic_vector(to_unsigned(174, 8)),
	3561 => std_logic_vector(to_unsigned(167, 8)),
	3562 => std_logic_vector(to_unsigned(165, 8)),
	3563 => std_logic_vector(to_unsigned(173, 8)),
	3564 => std_logic_vector(to_unsigned(165, 8)),
	3565 => std_logic_vector(to_unsigned(174, 8)),
	3566 => std_logic_vector(to_unsigned(165, 8)),
	3567 => std_logic_vector(to_unsigned(170, 8)),
	3568 => std_logic_vector(to_unsigned(168, 8)),
	3569 => std_logic_vector(to_unsigned(164, 8)),
	3570 => std_logic_vector(to_unsigned(174, 8)),
	3571 => std_logic_vector(to_unsigned(165, 8)),
	3572 => std_logic_vector(to_unsigned(176, 8)),
	3573 => std_logic_vector(to_unsigned(169, 8)),
	3574 => std_logic_vector(to_unsigned(164, 8)),
	3575 => std_logic_vector(to_unsigned(171, 8)),
	3576 => std_logic_vector(to_unsigned(173, 8)),
	3577 => std_logic_vector(to_unsigned(174, 8)),
	3578 => std_logic_vector(to_unsigned(172, 8)),
	3579 => std_logic_vector(to_unsigned(166, 8)),
	3580 => std_logic_vector(to_unsigned(164, 8)),
	3581 => std_logic_vector(to_unsigned(163, 8)),
	3582 => std_logic_vector(to_unsigned(175, 8)),
	3583 => std_logic_vector(to_unsigned(163, 8)),
	3584 => std_logic_vector(to_unsigned(176, 8)),
	3585 => std_logic_vector(to_unsigned(175, 8)),
	3586 => std_logic_vector(to_unsigned(175, 8)),
	3587 => std_logic_vector(to_unsigned(168, 8)),
	3588 => std_logic_vector(to_unsigned(169, 8)),
	3589 => std_logic_vector(to_unsigned(162, 8)),
	3590 => std_logic_vector(to_unsigned(176, 8)),
	3591 => std_logic_vector(to_unsigned(175, 8)),
	3592 => std_logic_vector(to_unsigned(167, 8)),
	3593 => std_logic_vector(to_unsigned(176, 8)),
	3594 => std_logic_vector(to_unsigned(176, 8)),
	3595 => std_logic_vector(to_unsigned(163, 8)),
	3596 => std_logic_vector(to_unsigned(168, 8)),
	3597 => std_logic_vector(to_unsigned(164, 8)),
	3598 => std_logic_vector(to_unsigned(170, 8)),
	3599 => std_logic_vector(to_unsigned(167, 8)),
	3600 => std_logic_vector(to_unsigned(172, 8)),
	3601 => std_logic_vector(to_unsigned(168, 8)),
	3602 => std_logic_vector(to_unsigned(166, 8)),
	3603 => std_logic_vector(to_unsigned(170, 8)),
	3604 => std_logic_vector(to_unsigned(170, 8)),
	3605 => std_logic_vector(to_unsigned(164, 8)),
	3606 => std_logic_vector(to_unsigned(174, 8)),
	3607 => std_logic_vector(to_unsigned(167, 8)),
	3608 => std_logic_vector(to_unsigned(167, 8)),
	3609 => std_logic_vector(to_unsigned(172, 8)),
	3610 => std_logic_vector(to_unsigned(167, 8)),
	3611 => std_logic_vector(to_unsigned(175, 8)),
	3612 => std_logic_vector(to_unsigned(175, 8)),
	3613 => std_logic_vector(to_unsigned(174, 8)),
	3614 => std_logic_vector(to_unsigned(176, 8)),
	3615 => std_logic_vector(to_unsigned(174, 8)),
	3616 => std_logic_vector(to_unsigned(165, 8)),
	3617 => std_logic_vector(to_unsigned(171, 8)),
	3618 => std_logic_vector(to_unsigned(167, 8)),
	3619 => std_logic_vector(to_unsigned(168, 8)),
	3620 => std_logic_vector(to_unsigned(174, 8)),
	3621 => std_logic_vector(to_unsigned(175, 8)),
	3622 => std_logic_vector(to_unsigned(163, 8)),
	3623 => std_logic_vector(to_unsigned(166, 8)),
	3624 => std_logic_vector(to_unsigned(170, 8)),
	3625 => std_logic_vector(to_unsigned(176, 8)),
	3626 => std_logic_vector(to_unsigned(174, 8)),
	3627 => std_logic_vector(to_unsigned(170, 8)),
	3628 => std_logic_vector(to_unsigned(166, 8)),
	3629 => std_logic_vector(to_unsigned(173, 8)),
	3630 => std_logic_vector(to_unsigned(169, 8)),
	3631 => std_logic_vector(to_unsigned(163, 8)),
	3632 => std_logic_vector(to_unsigned(165, 8)),
	3633 => std_logic_vector(to_unsigned(164, 8)),
	3634 => std_logic_vector(to_unsigned(167, 8)),
	3635 => std_logic_vector(to_unsigned(175, 8)),
	3636 => std_logic_vector(to_unsigned(166, 8)),
	3637 => std_logic_vector(to_unsigned(174, 8)),
	3638 => std_logic_vector(to_unsigned(168, 8)),
	3639 => std_logic_vector(to_unsigned(162, 8)),
	3640 => std_logic_vector(to_unsigned(163, 8)),
	3641 => std_logic_vector(to_unsigned(164, 8)),
	3642 => std_logic_vector(to_unsigned(174, 8)),
	3643 => std_logic_vector(to_unsigned(175, 8)),
	3644 => std_logic_vector(to_unsigned(173, 8)),
	3645 => std_logic_vector(to_unsigned(167, 8)),
	3646 => std_logic_vector(to_unsigned(173, 8)),
	3647 => std_logic_vector(to_unsigned(163, 8)),
	3648 => std_logic_vector(to_unsigned(166, 8)),
	3649 => std_logic_vector(to_unsigned(162, 8)),
	3650 => std_logic_vector(to_unsigned(171, 8)),
	3651 => std_logic_vector(to_unsigned(174, 8)),
	3652 => std_logic_vector(to_unsigned(169, 8)),
	3653 => std_logic_vector(to_unsigned(168, 8)),
	3654 => std_logic_vector(to_unsigned(172, 8)),
	3655 => std_logic_vector(to_unsigned(167, 8)),
	3656 => std_logic_vector(to_unsigned(171, 8)),
	3657 => std_logic_vector(to_unsigned(163, 8)),
	3658 => std_logic_vector(to_unsigned(174, 8)),
	3659 => std_logic_vector(to_unsigned(170, 8)),
	3660 => std_logic_vector(to_unsigned(176, 8)),
	3661 => std_logic_vector(to_unsigned(172, 8)),
	3662 => std_logic_vector(to_unsigned(167, 8)),
	3663 => std_logic_vector(to_unsigned(176, 8)),
	3664 => std_logic_vector(to_unsigned(173, 8)),
	3665 => std_logic_vector(to_unsigned(173, 8)),
	3666 => std_logic_vector(to_unsigned(175, 8)),
	3667 => std_logic_vector(to_unsigned(174, 8)),
	3668 => std_logic_vector(to_unsigned(166, 8)),
	3669 => std_logic_vector(to_unsigned(162, 8)),
	3670 => std_logic_vector(to_unsigned(162, 8)),
	3671 => std_logic_vector(to_unsigned(176, 8)),
	3672 => std_logic_vector(to_unsigned(170, 8)),
	3673 => std_logic_vector(to_unsigned(171, 8)),
	3674 => std_logic_vector(to_unsigned(163, 8)),
	3675 => std_logic_vector(to_unsigned(173, 8)),
	3676 => std_logic_vector(to_unsigned(164, 8)),
	3677 => std_logic_vector(to_unsigned(164, 8)),
	3678 => std_logic_vector(to_unsigned(162, 8)),
	3679 => std_logic_vector(to_unsigned(172, 8)),
	3680 => std_logic_vector(to_unsigned(167, 8)),
	3681 => std_logic_vector(to_unsigned(162, 8)),
	3682 => std_logic_vector(to_unsigned(172, 8)),
	3683 => std_logic_vector(to_unsigned(174, 8)),
	3684 => std_logic_vector(to_unsigned(170, 8)),
	3685 => std_logic_vector(to_unsigned(167, 8)),
	3686 => std_logic_vector(to_unsigned(168, 8)),
	3687 => std_logic_vector(to_unsigned(173, 8)),
	3688 => std_logic_vector(to_unsigned(163, 8)),
	3689 => std_logic_vector(to_unsigned(175, 8)),
	3690 => std_logic_vector(to_unsigned(163, 8)),
	3691 => std_logic_vector(to_unsigned(174, 8)),
	3692 => std_logic_vector(to_unsigned(174, 8)),
	3693 => std_logic_vector(to_unsigned(164, 8)),
	3694 => std_logic_vector(to_unsigned(173, 8)),
	3695 => std_logic_vector(to_unsigned(172, 8)),
	3696 => std_logic_vector(to_unsigned(175, 8)),
	3697 => std_logic_vector(to_unsigned(170, 8)),
	3698 => std_logic_vector(to_unsigned(172, 8)),
	3699 => std_logic_vector(to_unsigned(172, 8)),
	3700 => std_logic_vector(to_unsigned(175, 8)),
	3701 => std_logic_vector(to_unsigned(165, 8)),
	3702 => std_logic_vector(to_unsigned(163, 8)),
	3703 => std_logic_vector(to_unsigned(162, 8)),
	3704 => std_logic_vector(to_unsigned(174, 8)),
	3705 => std_logic_vector(to_unsigned(170, 8)),
	3706 => std_logic_vector(to_unsigned(163, 8)),
	3707 => std_logic_vector(to_unsigned(173, 8)),
	3708 => std_logic_vector(to_unsigned(173, 8)),
	3709 => std_logic_vector(to_unsigned(167, 8)),
	3710 => std_logic_vector(to_unsigned(163, 8)),
	3711 => std_logic_vector(to_unsigned(165, 8)),
	3712 => std_logic_vector(to_unsigned(169, 8)),
	3713 => std_logic_vector(to_unsigned(165, 8)),
	3714 => std_logic_vector(to_unsigned(176, 8)),
	3715 => std_logic_vector(to_unsigned(167, 8)),
	3716 => std_logic_vector(to_unsigned(173, 8)),
	3717 => std_logic_vector(to_unsigned(168, 8)),
	3718 => std_logic_vector(to_unsigned(172, 8)),
	3719 => std_logic_vector(to_unsigned(171, 8)),
	3720 => std_logic_vector(to_unsigned(164, 8)),
	3721 => std_logic_vector(to_unsigned(164, 8)),
	3722 => std_logic_vector(to_unsigned(175, 8)),
	3723 => std_logic_vector(to_unsigned(169, 8)),
	3724 => std_logic_vector(to_unsigned(167, 8)),
	3725 => std_logic_vector(to_unsigned(164, 8)),
	3726 => std_logic_vector(to_unsigned(162, 8)),
	3727 => std_logic_vector(to_unsigned(163, 8)),
	3728 => std_logic_vector(to_unsigned(169, 8)),
	3729 => std_logic_vector(to_unsigned(171, 8)),
	3730 => std_logic_vector(to_unsigned(171, 8)),
	3731 => std_logic_vector(to_unsigned(176, 8)),
	3732 => std_logic_vector(to_unsigned(174, 8)),
	3733 => std_logic_vector(to_unsigned(169, 8)),
	3734 => std_logic_vector(to_unsigned(170, 8)),
	3735 => std_logic_vector(to_unsigned(175, 8)),
	3736 => std_logic_vector(to_unsigned(169, 8)),
	3737 => std_logic_vector(to_unsigned(172, 8)),
	3738 => std_logic_vector(to_unsigned(171, 8)),
	3739 => std_logic_vector(to_unsigned(167, 8)),
	3740 => std_logic_vector(to_unsigned(170, 8)),
	3741 => std_logic_vector(to_unsigned(166, 8)),
	3742 => std_logic_vector(to_unsigned(165, 8)),
	3743 => std_logic_vector(to_unsigned(168, 8)),
	3744 => std_logic_vector(to_unsigned(171, 8)),
	3745 => std_logic_vector(to_unsigned(172, 8)),
	3746 => std_logic_vector(to_unsigned(165, 8)),
	3747 => std_logic_vector(to_unsigned(174, 8)),
	3748 => std_logic_vector(to_unsigned(174, 8)),
	3749 => std_logic_vector(to_unsigned(170, 8)),
	3750 => std_logic_vector(to_unsigned(163, 8)),
	3751 => std_logic_vector(to_unsigned(163, 8)),
	3752 => std_logic_vector(to_unsigned(173, 8)),
	3753 => std_logic_vector(to_unsigned(170, 8)),
	3754 => std_logic_vector(to_unsigned(175, 8)),
	3755 => std_logic_vector(to_unsigned(172, 8)),
	3756 => std_logic_vector(to_unsigned(169, 8)),
	3757 => std_logic_vector(to_unsigned(170, 8)),
	3758 => std_logic_vector(to_unsigned(174, 8)),
	3759 => std_logic_vector(to_unsigned(175, 8)),
	3760 => std_logic_vector(to_unsigned(171, 8)),
	3761 => std_logic_vector(to_unsigned(176, 8)),
	3762 => std_logic_vector(to_unsigned(163, 8)),
	3763 => std_logic_vector(to_unsigned(173, 8)),
	3764 => std_logic_vector(to_unsigned(175, 8)),
	3765 => std_logic_vector(to_unsigned(170, 8)),
	3766 => std_logic_vector(to_unsigned(169, 8)),
	3767 => std_logic_vector(to_unsigned(162, 8)),
	3768 => std_logic_vector(to_unsigned(171, 8)),
	3769 => std_logic_vector(to_unsigned(176, 8)),
	3770 => std_logic_vector(to_unsigned(175, 8)),
	3771 => std_logic_vector(to_unsigned(162, 8)),
	3772 => std_logic_vector(to_unsigned(169, 8)),
	3773 => std_logic_vector(to_unsigned(167, 8)),
	3774 => std_logic_vector(to_unsigned(164, 8)),
	3775 => std_logic_vector(to_unsigned(165, 8)),
	3776 => std_logic_vector(to_unsigned(172, 8)),
	3777 => std_logic_vector(to_unsigned(167, 8)),
	3778 => std_logic_vector(to_unsigned(174, 8)),
	3779 => std_logic_vector(to_unsigned(174, 8)),
	3780 => std_logic_vector(to_unsigned(176, 8)),
	3781 => std_logic_vector(to_unsigned(169, 8)),
	3782 => std_logic_vector(to_unsigned(168, 8)),
	3783 => std_logic_vector(to_unsigned(175, 8)),
	3784 => std_logic_vector(to_unsigned(176, 8)),
	3785 => std_logic_vector(to_unsigned(175, 8)),
	3786 => std_logic_vector(to_unsigned(174, 8)),
	3787 => std_logic_vector(to_unsigned(171, 8)),
	3788 => std_logic_vector(to_unsigned(176, 8)),
	3789 => std_logic_vector(to_unsigned(168, 8)),
	3790 => std_logic_vector(to_unsigned(172, 8)),
	3791 => std_logic_vector(to_unsigned(165, 8)),
	3792 => std_logic_vector(to_unsigned(163, 8)),
	3793 => std_logic_vector(to_unsigned(168, 8)),
	3794 => std_logic_vector(to_unsigned(162, 8)),
	3795 => std_logic_vector(to_unsigned(174, 8)),
	3796 => std_logic_vector(to_unsigned(166, 8)),
	3797 => std_logic_vector(to_unsigned(173, 8)),
	3798 => std_logic_vector(to_unsigned(174, 8)),
	3799 => std_logic_vector(to_unsigned(163, 8)),
	3800 => std_logic_vector(to_unsigned(175, 8)),
	3801 => std_logic_vector(to_unsigned(163, 8)),
	3802 => std_logic_vector(to_unsigned(175, 8)),
	3803 => std_logic_vector(to_unsigned(175, 8)),
	3804 => std_logic_vector(to_unsigned(166, 8)),
	3805 => std_logic_vector(to_unsigned(174, 8)),
	3806 => std_logic_vector(to_unsigned(175, 8)),
	3807 => std_logic_vector(to_unsigned(168, 8)),
	3808 => std_logic_vector(to_unsigned(167, 8)),
	3809 => std_logic_vector(to_unsigned(171, 8)),
	3810 => std_logic_vector(to_unsigned(165, 8)),
	3811 => std_logic_vector(to_unsigned(171, 8)),
	3812 => std_logic_vector(to_unsigned(167, 8)),
	3813 => std_logic_vector(to_unsigned(168, 8)),
	3814 => std_logic_vector(to_unsigned(163, 8)),
	3815 => std_logic_vector(to_unsigned(174, 8)),
	3816 => std_logic_vector(to_unsigned(176, 8)),
	3817 => std_logic_vector(to_unsigned(168, 8)),
	3818 => std_logic_vector(to_unsigned(162, 8)),
	3819 => std_logic_vector(to_unsigned(174, 8)),
	3820 => std_logic_vector(to_unsigned(164, 8)),
	3821 => std_logic_vector(to_unsigned(164, 8)),
	3822 => std_logic_vector(to_unsigned(176, 8)),
	3823 => std_logic_vector(to_unsigned(166, 8)),
	3824 => std_logic_vector(to_unsigned(171, 8)),
	3825 => std_logic_vector(to_unsigned(166, 8)),
	3826 => std_logic_vector(to_unsigned(170, 8)),
	3827 => std_logic_vector(to_unsigned(169, 8)),
	3828 => std_logic_vector(to_unsigned(176, 8)),
	3829 => std_logic_vector(to_unsigned(168, 8)),
	3830 => std_logic_vector(to_unsigned(170, 8)),
	3831 => std_logic_vector(to_unsigned(166, 8)),
	3832 => std_logic_vector(to_unsigned(169, 8)),
	3833 => std_logic_vector(to_unsigned(173, 8)),
	3834 => std_logic_vector(to_unsigned(174, 8)),
	3835 => std_logic_vector(to_unsigned(166, 8)),
	3836 => std_logic_vector(to_unsigned(170, 8)),
	3837 => std_logic_vector(to_unsigned(164, 8)),
	3838 => std_logic_vector(to_unsigned(165, 8)),
	3839 => std_logic_vector(to_unsigned(162, 8)),
	3840 => std_logic_vector(to_unsigned(172, 8)),
	3841 => std_logic_vector(to_unsigned(164, 8)),
	3842 => std_logic_vector(to_unsigned(168, 8)),
	3843 => std_logic_vector(to_unsigned(171, 8)),
	3844 => std_logic_vector(to_unsigned(169, 8)),
	3845 => std_logic_vector(to_unsigned(164, 8)),
	3846 => std_logic_vector(to_unsigned(167, 8)),
	3847 => std_logic_vector(to_unsigned(162, 8)),
	3848 => std_logic_vector(to_unsigned(165, 8)),
	3849 => std_logic_vector(to_unsigned(167, 8)),
	3850 => std_logic_vector(to_unsigned(168, 8)),
	3851 => std_logic_vector(to_unsigned(162, 8)),
	3852 => std_logic_vector(to_unsigned(164, 8)),
	3853 => std_logic_vector(to_unsigned(164, 8)),
	3854 => std_logic_vector(to_unsigned(175, 8)),
	3855 => std_logic_vector(to_unsigned(171, 8)),
	3856 => std_logic_vector(to_unsigned(168, 8)),
	3857 => std_logic_vector(to_unsigned(166, 8)),
	3858 => std_logic_vector(to_unsigned(174, 8)),
	3859 => std_logic_vector(to_unsigned(162, 8)),
	3860 => std_logic_vector(to_unsigned(170, 8)),
	3861 => std_logic_vector(to_unsigned(172, 8)),
	3862 => std_logic_vector(to_unsigned(171, 8)),
	3863 => std_logic_vector(to_unsigned(173, 8)),
	3864 => std_logic_vector(to_unsigned(170, 8)),
	3865 => std_logic_vector(to_unsigned(164, 8)),
	3866 => std_logic_vector(to_unsigned(169, 8)),
	3867 => std_logic_vector(to_unsigned(174, 8)),
	3868 => std_logic_vector(to_unsigned(165, 8)),
	3869 => std_logic_vector(to_unsigned(173, 8)),
	3870 => std_logic_vector(to_unsigned(162, 8)),
	3871 => std_logic_vector(to_unsigned(169, 8)),
	3872 => std_logic_vector(to_unsigned(167, 8)),
	3873 => std_logic_vector(to_unsigned(162, 8)),
	3874 => std_logic_vector(to_unsigned(167, 8)),
	3875 => std_logic_vector(to_unsigned(170, 8)),
	3876 => std_logic_vector(to_unsigned(176, 8)),
	3877 => std_logic_vector(to_unsigned(163, 8)),
	3878 => std_logic_vector(to_unsigned(169, 8)),
	3879 => std_logic_vector(to_unsigned(166, 8)),
	3880 => std_logic_vector(to_unsigned(162, 8)),
	3881 => std_logic_vector(to_unsigned(163, 8)),
	3882 => std_logic_vector(to_unsigned(171, 8)),
	3883 => std_logic_vector(to_unsigned(176, 8)),
	3884 => std_logic_vector(to_unsigned(165, 8)),
	3885 => std_logic_vector(to_unsigned(166, 8)),
	3886 => std_logic_vector(to_unsigned(168, 8)),
	3887 => std_logic_vector(to_unsigned(173, 8)),
	3888 => std_logic_vector(to_unsigned(162, 8)),
	3889 => std_logic_vector(to_unsigned(173, 8)),
	3890 => std_logic_vector(to_unsigned(175, 8)),
	3891 => std_logic_vector(to_unsigned(163, 8)),
	3892 => std_logic_vector(to_unsigned(164, 8)),
	3893 => std_logic_vector(to_unsigned(166, 8)),
	3894 => std_logic_vector(to_unsigned(164, 8)),
	3895 => std_logic_vector(to_unsigned(163, 8)),
	3896 => std_logic_vector(to_unsigned(164, 8)),
	3897 => std_logic_vector(to_unsigned(162, 8)),
	3898 => std_logic_vector(to_unsigned(169, 8)),
	3899 => std_logic_vector(to_unsigned(169, 8)),
	3900 => std_logic_vector(to_unsigned(164, 8)),
	3901 => std_logic_vector(to_unsigned(167, 8)),
	3902 => std_logic_vector(to_unsigned(173, 8)),
	3903 => std_logic_vector(to_unsigned(162, 8)),
	3904 => std_logic_vector(to_unsigned(168, 8)),
	3905 => std_logic_vector(to_unsigned(168, 8)),
	3906 => std_logic_vector(to_unsigned(170, 8)),
	3907 => std_logic_vector(to_unsigned(175, 8)),
	3908 => std_logic_vector(to_unsigned(164, 8)),
	3909 => std_logic_vector(to_unsigned(175, 8)),
	3910 => std_logic_vector(to_unsigned(171, 8)),
	3911 => std_logic_vector(to_unsigned(175, 8)),
	3912 => std_logic_vector(to_unsigned(170, 8)),
	3913 => std_logic_vector(to_unsigned(162, 8)),
	3914 => std_logic_vector(to_unsigned(170, 8)),
	3915 => std_logic_vector(to_unsigned(164, 8)),
	3916 => std_logic_vector(to_unsigned(164, 8)),
	3917 => std_logic_vector(to_unsigned(173, 8)),
	3918 => std_logic_vector(to_unsigned(176, 8)),
	3919 => std_logic_vector(to_unsigned(176, 8)),
	3920 => std_logic_vector(to_unsigned(169, 8)),
	3921 => std_logic_vector(to_unsigned(168, 8)),
	3922 => std_logic_vector(to_unsigned(162, 8)),
	3923 => std_logic_vector(to_unsigned(171, 8)),
	3924 => std_logic_vector(to_unsigned(163, 8)),
	3925 => std_logic_vector(to_unsigned(173, 8)),
	3926 => std_logic_vector(to_unsigned(169, 8)),
	3927 => std_logic_vector(to_unsigned(172, 8)),
	3928 => std_logic_vector(to_unsigned(162, 8)),
	3929 => std_logic_vector(to_unsigned(174, 8)),
	3930 => std_logic_vector(to_unsigned(166, 8)),
	3931 => std_logic_vector(to_unsigned(166, 8)),
	3932 => std_logic_vector(to_unsigned(170, 8)),
	3933 => std_logic_vector(to_unsigned(167, 8)),
	3934 => std_logic_vector(to_unsigned(171, 8)),
	3935 => std_logic_vector(to_unsigned(166, 8)),
	3936 => std_logic_vector(to_unsigned(171, 8)),
	3937 => std_logic_vector(to_unsigned(176, 8)),
	3938 => std_logic_vector(to_unsigned(165, 8)),
	3939 => std_logic_vector(to_unsigned(176, 8)),
	3940 => std_logic_vector(to_unsigned(167, 8)),
	3941 => std_logic_vector(to_unsigned(174, 8)),
	3942 => std_logic_vector(to_unsigned(176, 8)),
	3943 => std_logic_vector(to_unsigned(172, 8)),
	3944 => std_logic_vector(to_unsigned(164, 8)),
	3945 => std_logic_vector(to_unsigned(172, 8)),
	3946 => std_logic_vector(to_unsigned(170, 8)),
	3947 => std_logic_vector(to_unsigned(173, 8)),
	3948 => std_logic_vector(to_unsigned(175, 8)),
	3949 => std_logic_vector(to_unsigned(175, 8)),
	3950 => std_logic_vector(to_unsigned(171, 8)),
	3951 => std_logic_vector(to_unsigned(168, 8)),
	3952 => std_logic_vector(to_unsigned(168, 8)),
	3953 => std_logic_vector(to_unsigned(167, 8)),
	3954 => std_logic_vector(to_unsigned(173, 8)),
	3955 => std_logic_vector(to_unsigned(176, 8)),
	3956 => std_logic_vector(to_unsigned(164, 8)),
	3957 => std_logic_vector(to_unsigned(175, 8)),
	3958 => std_logic_vector(to_unsigned(166, 8)),
	3959 => std_logic_vector(to_unsigned(172, 8)),
	3960 => std_logic_vector(to_unsigned(171, 8)),
	3961 => std_logic_vector(to_unsigned(163, 8)),
	3962 => std_logic_vector(to_unsigned(165, 8)),
	3963 => std_logic_vector(to_unsigned(170, 8)),
	3964 => std_logic_vector(to_unsigned(164, 8)),
	3965 => std_logic_vector(to_unsigned(173, 8)),
	3966 => std_logic_vector(to_unsigned(166, 8)),
	3967 => std_logic_vector(to_unsigned(176, 8)),
	3968 => std_logic_vector(to_unsigned(164, 8)),
	3969 => std_logic_vector(to_unsigned(168, 8)),
	3970 => std_logic_vector(to_unsigned(173, 8)),
	3971 => std_logic_vector(to_unsigned(167, 8)),
	3972 => std_logic_vector(to_unsigned(176, 8)),
	3973 => std_logic_vector(to_unsigned(175, 8)),
	3974 => std_logic_vector(to_unsigned(164, 8)),
	3975 => std_logic_vector(to_unsigned(176, 8)),
	3976 => std_logic_vector(to_unsigned(170, 8)),
	3977 => std_logic_vector(to_unsigned(170, 8)),
	3978 => std_logic_vector(to_unsigned(175, 8)),
	3979 => std_logic_vector(to_unsigned(162, 8)),
	3980 => std_logic_vector(to_unsigned(167, 8)),
	3981 => std_logic_vector(to_unsigned(163, 8)),
	3982 => std_logic_vector(to_unsigned(176, 8)),
	3983 => std_logic_vector(to_unsigned(174, 8)),
	3984 => std_logic_vector(to_unsigned(171, 8)),
	3985 => std_logic_vector(to_unsigned(170, 8)),
	3986 => std_logic_vector(to_unsigned(163, 8)),
	3987 => std_logic_vector(to_unsigned(168, 8)),
	3988 => std_logic_vector(to_unsigned(173, 8)),
	3989 => std_logic_vector(to_unsigned(174, 8)),
	3990 => std_logic_vector(to_unsigned(170, 8)),
	3991 => std_logic_vector(to_unsigned(167, 8)),
	3992 => std_logic_vector(to_unsigned(176, 8)),
	3993 => std_logic_vector(to_unsigned(169, 8)),
	3994 => std_logic_vector(to_unsigned(172, 8)),
	3995 => std_logic_vector(to_unsigned(174, 8)),
	3996 => std_logic_vector(to_unsigned(162, 8)),
	3997 => std_logic_vector(to_unsigned(172, 8)),
	3998 => std_logic_vector(to_unsigned(175, 8)),
	3999 => std_logic_vector(to_unsigned(174, 8)),
	4000 => std_logic_vector(to_unsigned(165, 8)),
	4001 => std_logic_vector(to_unsigned(163, 8)),
	4002 => std_logic_vector(to_unsigned(176, 8)),
	4003 => std_logic_vector(to_unsigned(169, 8)),
	4004 => std_logic_vector(to_unsigned(170, 8)),
	4005 => std_logic_vector(to_unsigned(176, 8)),
	4006 => std_logic_vector(to_unsigned(168, 8)),
	4007 => std_logic_vector(to_unsigned(172, 8)),
	4008 => std_logic_vector(to_unsigned(171, 8)),
	4009 => std_logic_vector(to_unsigned(170, 8)),
	4010 => std_logic_vector(to_unsigned(163, 8)),
	4011 => std_logic_vector(to_unsigned(172, 8)),
	4012 => std_logic_vector(to_unsigned(174, 8)),
	4013 => std_logic_vector(to_unsigned(175, 8)),
	4014 => std_logic_vector(to_unsigned(170, 8)),
	4015 => std_logic_vector(to_unsigned(173, 8)),
	4016 => std_logic_vector(to_unsigned(173, 8)),
	4017 => std_logic_vector(to_unsigned(172, 8)),
	4018 => std_logic_vector(to_unsigned(171, 8)),
	4019 => std_logic_vector(to_unsigned(176, 8)),
	4020 => std_logic_vector(to_unsigned(169, 8)),
	4021 => std_logic_vector(to_unsigned(169, 8)),
	4022 => std_logic_vector(to_unsigned(173, 8)),
	4023 => std_logic_vector(to_unsigned(171, 8)),
	4024 => std_logic_vector(to_unsigned(176, 8)),
	4025 => std_logic_vector(to_unsigned(162, 8)),
	4026 => std_logic_vector(to_unsigned(173, 8)),
	4027 => std_logic_vector(to_unsigned(163, 8)),
	4028 => std_logic_vector(to_unsigned(166, 8)),
	4029 => std_logic_vector(to_unsigned(162, 8)),
	4030 => std_logic_vector(to_unsigned(166, 8)),
	4031 => std_logic_vector(to_unsigned(163, 8)),
	4032 => std_logic_vector(to_unsigned(172, 8)),
	4033 => std_logic_vector(to_unsigned(165, 8)),
	4034 => std_logic_vector(to_unsigned(174, 8)),
	4035 => std_logic_vector(to_unsigned(167, 8)),
	4036 => std_logic_vector(to_unsigned(174, 8)),
	4037 => std_logic_vector(to_unsigned(165, 8)),
	4038 => std_logic_vector(to_unsigned(175, 8)),
	4039 => std_logic_vector(to_unsigned(172, 8)),
	4040 => std_logic_vector(to_unsigned(176, 8)),
	4041 => std_logic_vector(to_unsigned(176, 8)),
	4042 => std_logic_vector(to_unsigned(170, 8)),
	4043 => std_logic_vector(to_unsigned(175, 8)),
	4044 => std_logic_vector(to_unsigned(163, 8)),
	4045 => std_logic_vector(to_unsigned(164, 8)),
	4046 => std_logic_vector(to_unsigned(174, 8)),
	4047 => std_logic_vector(to_unsigned(173, 8)),
	4048 => std_logic_vector(to_unsigned(168, 8)),
	4049 => std_logic_vector(to_unsigned(176, 8)),
	4050 => std_logic_vector(to_unsigned(166, 8)),
	4051 => std_logic_vector(to_unsigned(162, 8)),
	4052 => std_logic_vector(to_unsigned(170, 8)),
	4053 => std_logic_vector(to_unsigned(171, 8)),
	4054 => std_logic_vector(to_unsigned(168, 8)),
	4055 => std_logic_vector(to_unsigned(173, 8)),
	4056 => std_logic_vector(to_unsigned(176, 8)),
	4057 => std_logic_vector(to_unsigned(162, 8)),
	4058 => std_logic_vector(to_unsigned(174, 8)),
	4059 => std_logic_vector(to_unsigned(163, 8)),
	4060 => std_logic_vector(to_unsigned(163, 8)),
	4061 => std_logic_vector(to_unsigned(175, 8)),
	4062 => std_logic_vector(to_unsigned(169, 8)),
	4063 => std_logic_vector(to_unsigned(164, 8)),
	4064 => std_logic_vector(to_unsigned(176, 8)),
	4065 => std_logic_vector(to_unsigned(173, 8)),
	4066 => std_logic_vector(to_unsigned(168, 8)),
	4067 => std_logic_vector(to_unsigned(162, 8)),
	4068 => std_logic_vector(to_unsigned(162, 8)),
	4069 => std_logic_vector(to_unsigned(162, 8)),
	4070 => std_logic_vector(to_unsigned(171, 8)),
	4071 => std_logic_vector(to_unsigned(163, 8)),
	4072 => std_logic_vector(to_unsigned(169, 8)),
	4073 => std_logic_vector(to_unsigned(173, 8)),
	4074 => std_logic_vector(to_unsigned(168, 8)),
	4075 => std_logic_vector(to_unsigned(176, 8)),
	4076 => std_logic_vector(to_unsigned(176, 8)),
	4077 => std_logic_vector(to_unsigned(175, 8)),
	4078 => std_logic_vector(to_unsigned(162, 8)),
	4079 => std_logic_vector(to_unsigned(167, 8)),
	4080 => std_logic_vector(to_unsigned(162, 8)),
	4081 => std_logic_vector(to_unsigned(162, 8)),
	4082 => std_logic_vector(to_unsigned(165, 8)),
	4083 => std_logic_vector(to_unsigned(170, 8)),
	4084 => std_logic_vector(to_unsigned(163, 8)),
	4085 => std_logic_vector(to_unsigned(166, 8)),
	4086 => std_logic_vector(to_unsigned(166, 8)),
	4087 => std_logic_vector(to_unsigned(174, 8)),
	4088 => std_logic_vector(to_unsigned(174, 8)),
	4089 => std_logic_vector(to_unsigned(171, 8)),
	4090 => std_logic_vector(to_unsigned(169, 8)),
	4091 => std_logic_vector(to_unsigned(167, 8)),
	4092 => std_logic_vector(to_unsigned(172, 8)),
	4093 => std_logic_vector(to_unsigned(169, 8)),
	4094 => std_logic_vector(to_unsigned(169, 8)),
	4095 => std_logic_vector(to_unsigned(163, 8)),
	4096 => std_logic_vector(to_unsigned(176, 8)),
	4097 => std_logic_vector(to_unsigned(174, 8)),
	4098 => std_logic_vector(to_unsigned(162, 8)),
	4099 => std_logic_vector(to_unsigned(163, 8)),
	4100 => std_logic_vector(to_unsigned(167, 8)),
	4101 => std_logic_vector(to_unsigned(176, 8)),
	4102 => std_logic_vector(to_unsigned(168, 8)),
	4103 => std_logic_vector(to_unsigned(163, 8)),
	4104 => std_logic_vector(to_unsigned(170, 8)),
	4105 => std_logic_vector(to_unsigned(168, 8)),
	4106 => std_logic_vector(to_unsigned(175, 8)),
	4107 => std_logic_vector(to_unsigned(164, 8)),
	4108 => std_logic_vector(to_unsigned(176, 8)),
	4109 => std_logic_vector(to_unsigned(168, 8)),
	4110 => std_logic_vector(to_unsigned(174, 8)),
	4111 => std_logic_vector(to_unsigned(176, 8)),
	4112 => std_logic_vector(to_unsigned(172, 8)),
	4113 => std_logic_vector(to_unsigned(169, 8)),
	4114 => std_logic_vector(to_unsigned(169, 8)),
	4115 => std_logic_vector(to_unsigned(166, 8)),
	4116 => std_logic_vector(to_unsigned(162, 8)),
	4117 => std_logic_vector(to_unsigned(172, 8)),
	4118 => std_logic_vector(to_unsigned(173, 8)),
	4119 => std_logic_vector(to_unsigned(165, 8)),
	4120 => std_logic_vector(to_unsigned(168, 8)),
	4121 => std_logic_vector(to_unsigned(173, 8)),
	4122 => std_logic_vector(to_unsigned(174, 8)),
	4123 => std_logic_vector(to_unsigned(173, 8)),
	4124 => std_logic_vector(to_unsigned(176, 8)),
	4125 => std_logic_vector(to_unsigned(172, 8)),
	4126 => std_logic_vector(to_unsigned(175, 8)),
	4127 => std_logic_vector(to_unsigned(172, 8)),
	4128 => std_logic_vector(to_unsigned(164, 8)),
	4129 => std_logic_vector(to_unsigned(170, 8)),
	4130 => std_logic_vector(to_unsigned(173, 8)),
	4131 => std_logic_vector(to_unsigned(168, 8)),
	4132 => std_logic_vector(to_unsigned(164, 8)),
	4133 => std_logic_vector(to_unsigned(175, 8)),
	4134 => std_logic_vector(to_unsigned(164, 8)),
	4135 => std_logic_vector(to_unsigned(176, 8)),
	4136 => std_logic_vector(to_unsigned(173, 8)),
	4137 => std_logic_vector(to_unsigned(168, 8)),
	4138 => std_logic_vector(to_unsigned(165, 8)),
	4139 => std_logic_vector(to_unsigned(167, 8)),
	4140 => std_logic_vector(to_unsigned(176, 8)),
	4141 => std_logic_vector(to_unsigned(175, 8)),
	4142 => std_logic_vector(to_unsigned(164, 8)),
	4143 => std_logic_vector(to_unsigned(176, 8)),
	4144 => std_logic_vector(to_unsigned(163, 8)),
	4145 => std_logic_vector(to_unsigned(165, 8)),
	4146 => std_logic_vector(to_unsigned(163, 8)),
	4147 => std_logic_vector(to_unsigned(174, 8)),
	4148 => std_logic_vector(to_unsigned(175, 8)),
	4149 => std_logic_vector(to_unsigned(171, 8)),
	4150 => std_logic_vector(to_unsigned(164, 8)),
	4151 => std_logic_vector(to_unsigned(174, 8)),
	4152 => std_logic_vector(to_unsigned(171, 8)),
	4153 => std_logic_vector(to_unsigned(170, 8)),
	4154 => std_logic_vector(to_unsigned(168, 8)),
	4155 => std_logic_vector(to_unsigned(163, 8)),
	4156 => std_logic_vector(to_unsigned(175, 8)),
	4157 => std_logic_vector(to_unsigned(164, 8)),
	4158 => std_logic_vector(to_unsigned(167, 8)),
	4159 => std_logic_vector(to_unsigned(171, 8)),
	4160 => std_logic_vector(to_unsigned(162, 8)),
	4161 => std_logic_vector(to_unsigned(165, 8)),
	4162 => std_logic_vector(to_unsigned(168, 8)),
	4163 => std_logic_vector(to_unsigned(173, 8)),
	4164 => std_logic_vector(to_unsigned(163, 8)),
	4165 => std_logic_vector(to_unsigned(164, 8)),
	4166 => std_logic_vector(to_unsigned(172, 8)),
	4167 => std_logic_vector(to_unsigned(169, 8)),
	4168 => std_logic_vector(to_unsigned(175, 8)),
	4169 => std_logic_vector(to_unsigned(166, 8)),
	4170 => std_logic_vector(to_unsigned(175, 8)),
	4171 => std_logic_vector(to_unsigned(176, 8)),
	4172 => std_logic_vector(to_unsigned(164, 8)),
	4173 => std_logic_vector(to_unsigned(163, 8)),
	4174 => std_logic_vector(to_unsigned(168, 8)),
	4175 => std_logic_vector(to_unsigned(168, 8)),
	4176 => std_logic_vector(to_unsigned(176, 8)),
	4177 => std_logic_vector(to_unsigned(162, 8)),
	4178 => std_logic_vector(to_unsigned(170, 8)),
	4179 => std_logic_vector(to_unsigned(174, 8)),
	4180 => std_logic_vector(to_unsigned(170, 8)),
	4181 => std_logic_vector(to_unsigned(168, 8)),
	4182 => std_logic_vector(to_unsigned(168, 8)),
	4183 => std_logic_vector(to_unsigned(176, 8)),
	4184 => std_logic_vector(to_unsigned(166, 8)),
	4185 => std_logic_vector(to_unsigned(165, 8)),
	4186 => std_logic_vector(to_unsigned(169, 8)),
	4187 => std_logic_vector(to_unsigned(176, 8)),
	4188 => std_logic_vector(to_unsigned(171, 8)),
	4189 => std_logic_vector(to_unsigned(173, 8)),
	4190 => std_logic_vector(to_unsigned(168, 8)),
	others =>(others =>'0'));

component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_rst         : in  std_logic;
      i_start       : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector (7 downto 0)
      );
end component project_reti_logiche;


begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_rst      	=> tb_rst,
          i_start       => tb_start,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
          o_we 		=> mem_we,
          o_data    	=> mem_i_data
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;


MEM : process(tb_clk)
begin
    if tb_clk'event and tb_clk = '1' then
        if enable_wire = '1' then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
            end if;
        end if;
    end if;
end process;


test : process is
begin
    wait for 55 ns;
    -- wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    -- wait for c_CLOCK_PERIOD;
    -- wait for 100 ns;
    wait for 10 ns;
    tb_rst <= '0';
    -- wait for c_CLOCK_PERIOD;
    -- wait for 100 ns;
    tb_start <= '1';
    -- wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    -- wait for c_CLOCK_PERIOD;
    wait for 10 ns;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;

    assert RAM(4191) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4191)))) severity failure;
    assert RAM(4192) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4192)))) severity failure;
    assert RAM(4193) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4193)))) severity failure;
    assert RAM(4194) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4194)))) severity failure;
    assert RAM(4195) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4195)))) severity failure;
    assert RAM(4196) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4196)))) severity failure;
    assert RAM(4197) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4197)))) severity failure;
    assert RAM(4198) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4198)))) severity failure;
    assert RAM(4199) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4199)))) severity failure;
    assert RAM(4200) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4200)))) severity failure;
    assert RAM(4201) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4201)))) severity failure;
    assert RAM(4202) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4202)))) severity failure;
    assert RAM(4203) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4203)))) severity failure;
    assert RAM(4204) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4204)))) severity failure;
    assert RAM(4205) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4205)))) severity failure;
    assert RAM(4206) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4206)))) severity failure;
    assert RAM(4207) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4207)))) severity failure;
    assert RAM(4208) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4208)))) severity failure;
    assert RAM(4209) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4209)))) severity failure;
    assert RAM(4210) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4210)))) severity failure;
    assert RAM(4211) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4211)))) severity failure;
    assert RAM(4212) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4212)))) severity failure;
    assert RAM(4213) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4213)))) severity failure;
    assert RAM(4214) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4214)))) severity failure;
    assert RAM(4215) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4215)))) severity failure;
    assert RAM(4216) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4216)))) severity failure;
    assert RAM(4217) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4217)))) severity failure;
    assert RAM(4218) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4218)))) severity failure;
    assert RAM(4219) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4219)))) severity failure;
    assert RAM(4220) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4220)))) severity failure;
    assert RAM(4221) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4221)))) severity failure;
    assert RAM(4222) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4222)))) severity failure;
    assert RAM(4223) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4223)))) severity failure;
    assert RAM(4224) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4224)))) severity failure;
    assert RAM(4225) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4225)))) severity failure;
    assert RAM(4226) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4226)))) severity failure;
    assert RAM(4227) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4227)))) severity failure;
    assert RAM(4228) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4228)))) severity failure;
    assert RAM(4229) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4229)))) severity failure;
    assert RAM(4230) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4230)))) severity failure;
    assert RAM(4231) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4231)))) severity failure;
    assert RAM(4232) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4232)))) severity failure;
    assert RAM(4233) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4233)))) severity failure;
    assert RAM(4234) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4234)))) severity failure;
    assert RAM(4235) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4235)))) severity failure;
    assert RAM(4236) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4236)))) severity failure;
    assert RAM(4237) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4237)))) severity failure;
    assert RAM(4238) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4238)))) severity failure;
    assert RAM(4239) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4239)))) severity failure;
    assert RAM(4240) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4240)))) severity failure;
    assert RAM(4241) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4241)))) severity failure;
    assert RAM(4242) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4242)))) severity failure;
    assert RAM(4243) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4243)))) severity failure;
    assert RAM(4244) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4244)))) severity failure;
    assert RAM(4245) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4245)))) severity failure;
    assert RAM(4246) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4246)))) severity failure;
    assert RAM(4247) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4247)))) severity failure;
    assert RAM(4248) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4248)))) severity failure;
    assert RAM(4249) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4249)))) severity failure;
    assert RAM(4250) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4250)))) severity failure;
    assert RAM(4251) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4251)))) severity failure;
    assert RAM(4252) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4252)))) severity failure;
    assert RAM(4253) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4253)))) severity failure;
    assert RAM(4254) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4254)))) severity failure;
    assert RAM(4255) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4255)))) severity failure;
    assert RAM(4256) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4256)))) severity failure;
    assert RAM(4257) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4257)))) severity failure;
    assert RAM(4258) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4258)))) severity failure;
    assert RAM(4259) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4259)))) severity failure;
    assert RAM(4260) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4260)))) severity failure;
    assert RAM(4261) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4261)))) severity failure;
    assert RAM(4262) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4262)))) severity failure;
    assert RAM(4263) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4263)))) severity failure;
    assert RAM(4264) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4264)))) severity failure;
    assert RAM(4265) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4265)))) severity failure;
    assert RAM(4266) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4266)))) severity failure;
    assert RAM(4267) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4267)))) severity failure;
    assert RAM(4268) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4268)))) severity failure;
    assert RAM(4269) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4269)))) severity failure;
    assert RAM(4270) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4270)))) severity failure;
    assert RAM(4271) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4271)))) severity failure;
    assert RAM(4272) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4272)))) severity failure;
    assert RAM(4273) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4273)))) severity failure;
    assert RAM(4274) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4274)))) severity failure;
    assert RAM(4275) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4275)))) severity failure;
    assert RAM(4276) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4276)))) severity failure;
    assert RAM(4277) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4277)))) severity failure;
    assert RAM(4278) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4278)))) severity failure;
    assert RAM(4279) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4279)))) severity failure;
    assert RAM(4280) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4280)))) severity failure;
    assert RAM(4281) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4281)))) severity failure;
    assert RAM(4282) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4282)))) severity failure;
    assert RAM(4283) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4283)))) severity failure;
    assert RAM(4284) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4284)))) severity failure;
    assert RAM(4285) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4285)))) severity failure;
    assert RAM(4286) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4286)))) severity failure;
    assert RAM(4287) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4287)))) severity failure;
    assert RAM(4288) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4288)))) severity failure;
    assert RAM(4289) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4289)))) severity failure;
    assert RAM(4290) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4290)))) severity failure;
    assert RAM(4291) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4291)))) severity failure;
    assert RAM(4292) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4292)))) severity failure;
    assert RAM(4293) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4293)))) severity failure;
    assert RAM(4294) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4294)))) severity failure;
    assert RAM(4295) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4295)))) severity failure;
    assert RAM(4296) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4296)))) severity failure;
    assert RAM(4297) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4297)))) severity failure;
    assert RAM(4298) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4298)))) severity failure;
    assert RAM(4299) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4299)))) severity failure;
    assert RAM(4300) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4300)))) severity failure;
    assert RAM(4301) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4301)))) severity failure;
    assert RAM(4302) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4302)))) severity failure;
    assert RAM(4303) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4303)))) severity failure;
    assert RAM(4304) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4304)))) severity failure;
    assert RAM(4305) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4305)))) severity failure;
    assert RAM(4306) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4306)))) severity failure;
    assert RAM(4307) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4307)))) severity failure;
    assert RAM(4308) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4308)))) severity failure;
    assert RAM(4309) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4309)))) severity failure;
    assert RAM(4310) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4310)))) severity failure;
    assert RAM(4311) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4311)))) severity failure;
    assert RAM(4312) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4312)))) severity failure;
    assert RAM(4313) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4313)))) severity failure;
    assert RAM(4314) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4314)))) severity failure;
    assert RAM(4315) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4315)))) severity failure;
    assert RAM(4316) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4316)))) severity failure;
    assert RAM(4317) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4317)))) severity failure;
    assert RAM(4318) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4318)))) severity failure;
    assert RAM(4319) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4319)))) severity failure;
    assert RAM(4320) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4320)))) severity failure;
    assert RAM(4321) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4321)))) severity failure;
    assert RAM(4322) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4322)))) severity failure;
    assert RAM(4323) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4323)))) severity failure;
    assert RAM(4324) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4324)))) severity failure;
    assert RAM(4325) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4325)))) severity failure;
    assert RAM(4326) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4326)))) severity failure;
    assert RAM(4327) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4327)))) severity failure;
    assert RAM(4328) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4328)))) severity failure;
    assert RAM(4329) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4329)))) severity failure;
    assert RAM(4330) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4330)))) severity failure;
    assert RAM(4331) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4331)))) severity failure;
    assert RAM(4332) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4332)))) severity failure;
    assert RAM(4333) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4333)))) severity failure;
    assert RAM(4334) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4334)))) severity failure;
    assert RAM(4335) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4335)))) severity failure;
    assert RAM(4336) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4336)))) severity failure;
    assert RAM(4337) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4337)))) severity failure;
    assert RAM(4338) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4338)))) severity failure;
    assert RAM(4339) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4339)))) severity failure;
    assert RAM(4340) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4340)))) severity failure;
    assert RAM(4341) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4341)))) severity failure;
    assert RAM(4342) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4342)))) severity failure;
    assert RAM(4343) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4343)))) severity failure;
    assert RAM(4344) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4344)))) severity failure;
    assert RAM(4345) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4345)))) severity failure;
    assert RAM(4346) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4346)))) severity failure;
    assert RAM(4347) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4347)))) severity failure;
    assert RAM(4348) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4348)))) severity failure;
    assert RAM(4349) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4349)))) severity failure;
    assert RAM(4350) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4350)))) severity failure;
    assert RAM(4351) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4351)))) severity failure;
    assert RAM(4352) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4352)))) severity failure;
    assert RAM(4353) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4353)))) severity failure;
    assert RAM(4354) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4354)))) severity failure;
    assert RAM(4355) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4355)))) severity failure;
    assert RAM(4356) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4356)))) severity failure;
    assert RAM(4357) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4357)))) severity failure;
    assert RAM(4358) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4358)))) severity failure;
    assert RAM(4359) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4359)))) severity failure;
    assert RAM(4360) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4360)))) severity failure;
    assert RAM(4361) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4361)))) severity failure;
    assert RAM(4362) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4362)))) severity failure;
    assert RAM(4363) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4363)))) severity failure;
    assert RAM(4364) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4364)))) severity failure;
    assert RAM(4365) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4365)))) severity failure;
    assert RAM(4366) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4366)))) severity failure;
    assert RAM(4367) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4367)))) severity failure;
    assert RAM(4368) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4368)))) severity failure;
    assert RAM(4369) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4369)))) severity failure;
    assert RAM(4370) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4370)))) severity failure;
    assert RAM(4371) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4371)))) severity failure;
    assert RAM(4372) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4372)))) severity failure;
    assert RAM(4373) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4373)))) severity failure;
    assert RAM(4374) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4374)))) severity failure;
    assert RAM(4375) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4375)))) severity failure;
    assert RAM(4376) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4376)))) severity failure;
    assert RAM(4377) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4377)))) severity failure;
    assert RAM(4378) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4378)))) severity failure;
    assert RAM(4379) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4379)))) severity failure;
    assert RAM(4380) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4380)))) severity failure;
    assert RAM(4381) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4381)))) severity failure;
    assert RAM(4382) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4382)))) severity failure;
    assert RAM(4383) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4383)))) severity failure;
    assert RAM(4384) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4384)))) severity failure;
    assert RAM(4385) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4385)))) severity failure;
    assert RAM(4386) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4386)))) severity failure;
    assert RAM(4387) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4387)))) severity failure;
    assert RAM(4388) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4388)))) severity failure;
    assert RAM(4389) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4389)))) severity failure;
    assert RAM(4390) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4390)))) severity failure;
    assert RAM(4391) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4391)))) severity failure;
    assert RAM(4392) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4392)))) severity failure;
    assert RAM(4393) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4393)))) severity failure;
    assert RAM(4394) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4394)))) severity failure;
    assert RAM(4395) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4395)))) severity failure;
    assert RAM(4396) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4396)))) severity failure;
    assert RAM(4397) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4397)))) severity failure;
    assert RAM(4398) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4398)))) severity failure;
    assert RAM(4399) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4399)))) severity failure;
    assert RAM(4400) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4400)))) severity failure;
    assert RAM(4401) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4401)))) severity failure;
    assert RAM(4402) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4402)))) severity failure;
    assert RAM(4403) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4403)))) severity failure;
    assert RAM(4404) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4404)))) severity failure;
    assert RAM(4405) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4405)))) severity failure;
    assert RAM(4406) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4406)))) severity failure;
    assert RAM(4407) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4407)))) severity failure;
    assert RAM(4408) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4408)))) severity failure;
    assert RAM(4409) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4409)))) severity failure;
    assert RAM(4410) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4410)))) severity failure;
    assert RAM(4411) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4411)))) severity failure;
    assert RAM(4412) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4412)))) severity failure;
    assert RAM(4413) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4413)))) severity failure;
    assert RAM(4414) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4414)))) severity failure;
    assert RAM(4415) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4415)))) severity failure;
    assert RAM(4416) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4416)))) severity failure;
    assert RAM(4417) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4417)))) severity failure;
    assert RAM(4418) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4418)))) severity failure;
    assert RAM(4419) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4419)))) severity failure;
    assert RAM(4420) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4420)))) severity failure;
    assert RAM(4421) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4421)))) severity failure;
    assert RAM(4422) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4422)))) severity failure;
    assert RAM(4423) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4423)))) severity failure;
    assert RAM(4424) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4424)))) severity failure;
    assert RAM(4425) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4425)))) severity failure;
    assert RAM(4426) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4426)))) severity failure;
    assert RAM(4427) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4427)))) severity failure;
    assert RAM(4428) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4428)))) severity failure;
    assert RAM(4429) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4429)))) severity failure;
    assert RAM(4430) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4430)))) severity failure;
    assert RAM(4431) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4431)))) severity failure;
    assert RAM(4432) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4432)))) severity failure;
    assert RAM(4433) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4433)))) severity failure;
    assert RAM(4434) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4434)))) severity failure;
    assert RAM(4435) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4435)))) severity failure;
    assert RAM(4436) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4436)))) severity failure;
    assert RAM(4437) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4437)))) severity failure;
    assert RAM(4438) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4438)))) severity failure;
    assert RAM(4439) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4439)))) severity failure;
    assert RAM(4440) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4440)))) severity failure;
    assert RAM(4441) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4441)))) severity failure;
    assert RAM(4442) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4442)))) severity failure;
    assert RAM(4443) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4443)))) severity failure;
    assert RAM(4444) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4444)))) severity failure;
    assert RAM(4445) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4445)))) severity failure;
    assert RAM(4446) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4446)))) severity failure;
    assert RAM(4447) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4447)))) severity failure;
    assert RAM(4448) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4448)))) severity failure;
    assert RAM(4449) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4449)))) severity failure;
    assert RAM(4450) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4450)))) severity failure;
    assert RAM(4451) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4451)))) severity failure;
    assert RAM(4452) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4452)))) severity failure;
    assert RAM(4453) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4453)))) severity failure;
    assert RAM(4454) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4454)))) severity failure;
    assert RAM(4455) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4455)))) severity failure;
    assert RAM(4456) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4456)))) severity failure;
    assert RAM(4457) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4457)))) severity failure;
    assert RAM(4458) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4458)))) severity failure;
    assert RAM(4459) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4459)))) severity failure;
    assert RAM(4460) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4460)))) severity failure;
    assert RAM(4461) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4461)))) severity failure;
    assert RAM(4462) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4462)))) severity failure;
    assert RAM(4463) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4463)))) severity failure;
    assert RAM(4464) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4464)))) severity failure;
    assert RAM(4465) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4465)))) severity failure;
    assert RAM(4466) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4466)))) severity failure;
    assert RAM(4467) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4467)))) severity failure;
    assert RAM(4468) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4468)))) severity failure;
    assert RAM(4469) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4469)))) severity failure;
    assert RAM(4470) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4470)))) severity failure;
    assert RAM(4471) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4471)))) severity failure;
    assert RAM(4472) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4472)))) severity failure;
    assert RAM(4473) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4473)))) severity failure;
    assert RAM(4474) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4474)))) severity failure;
    assert RAM(4475) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4475)))) severity failure;
    assert RAM(4476) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4476)))) severity failure;
    assert RAM(4477) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4477)))) severity failure;
    assert RAM(4478) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4478)))) severity failure;
    assert RAM(4479) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4479)))) severity failure;
    assert RAM(4480) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4480)))) severity failure;
    assert RAM(4481) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4481)))) severity failure;
    assert RAM(4482) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4482)))) severity failure;
    assert RAM(4483) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4483)))) severity failure;
    assert RAM(4484) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4484)))) severity failure;
    assert RAM(4485) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4485)))) severity failure;
    assert RAM(4486) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4486)))) severity failure;
    assert RAM(4487) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4487)))) severity failure;
    assert RAM(4488) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4488)))) severity failure;
    assert RAM(4489) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4489)))) severity failure;
    assert RAM(4490) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4490)))) severity failure;
    assert RAM(4491) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4491)))) severity failure;
    assert RAM(4492) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4492)))) severity failure;
    assert RAM(4493) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4493)))) severity failure;
    assert RAM(4494) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4494)))) severity failure;
    assert RAM(4495) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4495)))) severity failure;
    assert RAM(4496) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4496)))) severity failure;
    assert RAM(4497) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4497)))) severity failure;
    assert RAM(4498) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4498)))) severity failure;
    assert RAM(4499) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4499)))) severity failure;
    assert RAM(4500) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4500)))) severity failure;
    assert RAM(4501) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4501)))) severity failure;
    assert RAM(4502) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4502)))) severity failure;
    assert RAM(4503) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4503)))) severity failure;
    assert RAM(4504) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4504)))) severity failure;
    assert RAM(4505) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4505)))) severity failure;
    assert RAM(4506) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4506)))) severity failure;
    assert RAM(4507) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4507)))) severity failure;
    assert RAM(4508) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4508)))) severity failure;
    assert RAM(4509) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4509)))) severity failure;
    assert RAM(4510) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4510)))) severity failure;
    assert RAM(4511) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4511)))) severity failure;
    assert RAM(4512) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4512)))) severity failure;
    assert RAM(4513) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4513)))) severity failure;
    assert RAM(4514) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4514)))) severity failure;
    assert RAM(4515) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4515)))) severity failure;
    assert RAM(4516) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4516)))) severity failure;
    assert RAM(4517) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4517)))) severity failure;
    assert RAM(4518) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4518)))) severity failure;
    assert RAM(4519) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4519)))) severity failure;
    assert RAM(4520) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4520)))) severity failure;
    assert RAM(4521) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4521)))) severity failure;
    assert RAM(4522) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4522)))) severity failure;
    assert RAM(4523) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4523)))) severity failure;
    assert RAM(4524) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4524)))) severity failure;
    assert RAM(4525) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4525)))) severity failure;
    assert RAM(4526) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4526)))) severity failure;
    assert RAM(4527) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4527)))) severity failure;
    assert RAM(4528) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4528)))) severity failure;
    assert RAM(4529) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4529)))) severity failure;
    assert RAM(4530) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4530)))) severity failure;
    assert RAM(4531) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4531)))) severity failure;
    assert RAM(4532) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4532)))) severity failure;
    assert RAM(4533) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4533)))) severity failure;
    assert RAM(4534) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4534)))) severity failure;
    assert RAM(4535) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4535)))) severity failure;
    assert RAM(4536) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4536)))) severity failure;
    assert RAM(4537) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4537)))) severity failure;
    assert RAM(4538) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4538)))) severity failure;
    assert RAM(4539) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4539)))) severity failure;
    assert RAM(4540) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4540)))) severity failure;
    assert RAM(4541) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4541)))) severity failure;
    assert RAM(4542) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4542)))) severity failure;
    assert RAM(4543) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4543)))) severity failure;
    assert RAM(4544) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4544)))) severity failure;
    assert RAM(4545) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4545)))) severity failure;
    assert RAM(4546) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4546)))) severity failure;
    assert RAM(4547) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4547)))) severity failure;
    assert RAM(4548) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4548)))) severity failure;
    assert RAM(4549) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4549)))) severity failure;
    assert RAM(4550) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4550)))) severity failure;
    assert RAM(4551) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4551)))) severity failure;
    assert RAM(4552) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4552)))) severity failure;
    assert RAM(4553) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4553)))) severity failure;
    assert RAM(4554) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4554)))) severity failure;
    assert RAM(4555) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4555)))) severity failure;
    assert RAM(4556) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4556)))) severity failure;
    assert RAM(4557) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4557)))) severity failure;
    assert RAM(4558) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4558)))) severity failure;
    assert RAM(4559) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4559)))) severity failure;
    assert RAM(4560) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4560)))) severity failure;
    assert RAM(4561) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4561)))) severity failure;
    assert RAM(4562) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4562)))) severity failure;
    assert RAM(4563) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4563)))) severity failure;
    assert RAM(4564) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4564)))) severity failure;
    assert RAM(4565) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4565)))) severity failure;
    assert RAM(4566) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4566)))) severity failure;
    assert RAM(4567) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4567)))) severity failure;
    assert RAM(4568) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4568)))) severity failure;
    assert RAM(4569) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4569)))) severity failure;
    assert RAM(4570) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4570)))) severity failure;
    assert RAM(4571) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4571)))) severity failure;
    assert RAM(4572) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4572)))) severity failure;
    assert RAM(4573) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4573)))) severity failure;
    assert RAM(4574) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4574)))) severity failure;
    assert RAM(4575) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4575)))) severity failure;
    assert RAM(4576) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4576)))) severity failure;
    assert RAM(4577) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4577)))) severity failure;
    assert RAM(4578) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4578)))) severity failure;
    assert RAM(4579) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4579)))) severity failure;
    assert RAM(4580) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4580)))) severity failure;
    assert RAM(4581) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4581)))) severity failure;
    assert RAM(4582) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4582)))) severity failure;
    assert RAM(4583) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4583)))) severity failure;
    assert RAM(4584) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4584)))) severity failure;
    assert RAM(4585) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4585)))) severity failure;
    assert RAM(4586) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4586)))) severity failure;
    assert RAM(4587) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4587)))) severity failure;
    assert RAM(4588) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4588)))) severity failure;
    assert RAM(4589) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4589)))) severity failure;
    assert RAM(4590) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4590)))) severity failure;
    assert RAM(4591) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4591)))) severity failure;
    assert RAM(4592) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4592)))) severity failure;
    assert RAM(4593) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4593)))) severity failure;
    assert RAM(4594) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4594)))) severity failure;
    assert RAM(4595) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4595)))) severity failure;
    assert RAM(4596) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4596)))) severity failure;
    assert RAM(4597) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4597)))) severity failure;
    assert RAM(4598) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4598)))) severity failure;
    assert RAM(4599) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4599)))) severity failure;
    assert RAM(4600) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4600)))) severity failure;
    assert RAM(4601) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4601)))) severity failure;
    assert RAM(4602) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4602)))) severity failure;
    assert RAM(4603) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4603)))) severity failure;
    assert RAM(4604) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4604)))) severity failure;
    assert RAM(4605) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4605)))) severity failure;
    assert RAM(4606) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4606)))) severity failure;
    assert RAM(4607) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4607)))) severity failure;
    assert RAM(4608) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4608)))) severity failure;
    assert RAM(4609) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4609)))) severity failure;
    assert RAM(4610) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4610)))) severity failure;
    assert RAM(4611) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4611)))) severity failure;
    assert RAM(4612) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4612)))) severity failure;
    assert RAM(4613) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4613)))) severity failure;
    assert RAM(4614) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4614)))) severity failure;
    assert RAM(4615) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4615)))) severity failure;
    assert RAM(4616) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4616)))) severity failure;
    assert RAM(4617) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4617)))) severity failure;
    assert RAM(4618) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4618)))) severity failure;
    assert RAM(4619) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4619)))) severity failure;
    assert RAM(4620) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4620)))) severity failure;
    assert RAM(4621) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4621)))) severity failure;
    assert RAM(4622) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4622)))) severity failure;
    assert RAM(4623) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4623)))) severity failure;
    assert RAM(4624) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4624)))) severity failure;
    assert RAM(4625) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4625)))) severity failure;
    assert RAM(4626) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4626)))) severity failure;
    assert RAM(4627) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4627)))) severity failure;
    assert RAM(4628) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4628)))) severity failure;
    assert RAM(4629) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4629)))) severity failure;
    assert RAM(4630) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4630)))) severity failure;
    assert RAM(4631) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4631)))) severity failure;
    assert RAM(4632) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4632)))) severity failure;
    assert RAM(4633) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4633)))) severity failure;
    assert RAM(4634) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4634)))) severity failure;
    assert RAM(4635) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4635)))) severity failure;
    assert RAM(4636) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4636)))) severity failure;
    assert RAM(4637) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4637)))) severity failure;
    assert RAM(4638) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4638)))) severity failure;
    assert RAM(4639) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4639)))) severity failure;
    assert RAM(4640) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4640)))) severity failure;
    assert RAM(4641) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4641)))) severity failure;
    assert RAM(4642) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4642)))) severity failure;
    assert RAM(4643) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4643)))) severity failure;
    assert RAM(4644) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4644)))) severity failure;
    assert RAM(4645) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4645)))) severity failure;
    assert RAM(4646) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4646)))) severity failure;
    assert RAM(4647) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4647)))) severity failure;
    assert RAM(4648) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4648)))) severity failure;
    assert RAM(4649) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4649)))) severity failure;
    assert RAM(4650) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4650)))) severity failure;
    assert RAM(4651) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4651)))) severity failure;
    assert RAM(4652) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4652)))) severity failure;
    assert RAM(4653) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4653)))) severity failure;
    assert RAM(4654) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4654)))) severity failure;
    assert RAM(4655) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4655)))) severity failure;
    assert RAM(4656) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4656)))) severity failure;
    assert RAM(4657) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4657)))) severity failure;
    assert RAM(4658) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4658)))) severity failure;
    assert RAM(4659) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4659)))) severity failure;
    assert RAM(4660) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4660)))) severity failure;
    assert RAM(4661) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4661)))) severity failure;
    assert RAM(4662) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4662)))) severity failure;
    assert RAM(4663) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4663)))) severity failure;
    assert RAM(4664) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4664)))) severity failure;
    assert RAM(4665) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4665)))) severity failure;
    assert RAM(4666) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4666)))) severity failure;
    assert RAM(4667) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4667)))) severity failure;
    assert RAM(4668) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4668)))) severity failure;
    assert RAM(4669) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4669)))) severity failure;
    assert RAM(4670) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4670)))) severity failure;
    assert RAM(4671) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4671)))) severity failure;
    assert RAM(4672) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4672)))) severity failure;
    assert RAM(4673) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4673)))) severity failure;
    assert RAM(4674) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4674)))) severity failure;
    assert RAM(4675) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4675)))) severity failure;
    assert RAM(4676) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4676)))) severity failure;
    assert RAM(4677) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4677)))) severity failure;
    assert RAM(4678) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4678)))) severity failure;
    assert RAM(4679) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4679)))) severity failure;
    assert RAM(4680) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4680)))) severity failure;
    assert RAM(4681) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4681)))) severity failure;
    assert RAM(4682) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4682)))) severity failure;
    assert RAM(4683) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4683)))) severity failure;
    assert RAM(4684) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4684)))) severity failure;
    assert RAM(4685) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4685)))) severity failure;
    assert RAM(4686) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4686)))) severity failure;
    assert RAM(4687) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4687)))) severity failure;
    assert RAM(4688) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4688)))) severity failure;
    assert RAM(4689) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4689)))) severity failure;
    assert RAM(4690) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4690)))) severity failure;
    assert RAM(4691) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4691)))) severity failure;
    assert RAM(4692) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4692)))) severity failure;
    assert RAM(4693) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4693)))) severity failure;
    assert RAM(4694) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4694)))) severity failure;
    assert RAM(4695) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4695)))) severity failure;
    assert RAM(4696) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4696)))) severity failure;
    assert RAM(4697) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4697)))) severity failure;
    assert RAM(4698) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4698)))) severity failure;
    assert RAM(4699) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4699)))) severity failure;
    assert RAM(4700) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4700)))) severity failure;
    assert RAM(4701) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4701)))) severity failure;
    assert RAM(4702) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4702)))) severity failure;
    assert RAM(4703) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4703)))) severity failure;
    assert RAM(4704) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4704)))) severity failure;
    assert RAM(4705) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4705)))) severity failure;
    assert RAM(4706) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4706)))) severity failure;
    assert RAM(4707) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4707)))) severity failure;
    assert RAM(4708) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4708)))) severity failure;
    assert RAM(4709) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4709)))) severity failure;
    assert RAM(4710) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4710)))) severity failure;
    assert RAM(4711) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4711)))) severity failure;
    assert RAM(4712) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4712)))) severity failure;
    assert RAM(4713) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4713)))) severity failure;
    assert RAM(4714) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4714)))) severity failure;
    assert RAM(4715) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4715)))) severity failure;
    assert RAM(4716) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4716)))) severity failure;
    assert RAM(4717) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4717)))) severity failure;
    assert RAM(4718) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4718)))) severity failure;
    assert RAM(4719) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4719)))) severity failure;
    assert RAM(4720) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4720)))) severity failure;
    assert RAM(4721) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4721)))) severity failure;
    assert RAM(4722) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4722)))) severity failure;
    assert RAM(4723) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4723)))) severity failure;
    assert RAM(4724) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4724)))) severity failure;
    assert RAM(4725) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4725)))) severity failure;
    assert RAM(4726) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4726)))) severity failure;
    assert RAM(4727) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4727)))) severity failure;
    assert RAM(4728) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4728)))) severity failure;
    assert RAM(4729) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4729)))) severity failure;
    assert RAM(4730) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4730)))) severity failure;
    assert RAM(4731) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4731)))) severity failure;
    assert RAM(4732) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4732)))) severity failure;
    assert RAM(4733) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4733)))) severity failure;
    assert RAM(4734) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4734)))) severity failure;
    assert RAM(4735) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4735)))) severity failure;
    assert RAM(4736) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4736)))) severity failure;
    assert RAM(4737) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4737)))) severity failure;
    assert RAM(4738) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4738)))) severity failure;
    assert RAM(4739) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4739)))) severity failure;
    assert RAM(4740) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4740)))) severity failure;
    assert RAM(4741) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4741)))) severity failure;
    assert RAM(4742) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4742)))) severity failure;
    assert RAM(4743) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4743)))) severity failure;
    assert RAM(4744) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4744)))) severity failure;
    assert RAM(4745) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4745)))) severity failure;
    assert RAM(4746) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4746)))) severity failure;
    assert RAM(4747) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4747)))) severity failure;
    assert RAM(4748) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4748)))) severity failure;
    assert RAM(4749) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4749)))) severity failure;
    assert RAM(4750) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4750)))) severity failure;
    assert RAM(4751) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4751)))) severity failure;
    assert RAM(4752) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4752)))) severity failure;
    assert RAM(4753) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4753)))) severity failure;
    assert RAM(4754) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4754)))) severity failure;
    assert RAM(4755) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4755)))) severity failure;
    assert RAM(4756) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4756)))) severity failure;
    assert RAM(4757) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4757)))) severity failure;
    assert RAM(4758) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4758)))) severity failure;
    assert RAM(4759) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4759)))) severity failure;
    assert RAM(4760) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4760)))) severity failure;
    assert RAM(4761) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4761)))) severity failure;
    assert RAM(4762) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4762)))) severity failure;
    assert RAM(4763) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4763)))) severity failure;
    assert RAM(4764) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4764)))) severity failure;
    assert RAM(4765) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4765)))) severity failure;
    assert RAM(4766) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4766)))) severity failure;
    assert RAM(4767) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4767)))) severity failure;
    assert RAM(4768) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4768)))) severity failure;
    assert RAM(4769) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4769)))) severity failure;
    assert RAM(4770) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4770)))) severity failure;
    assert RAM(4771) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4771)))) severity failure;
    assert RAM(4772) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4772)))) severity failure;
    assert RAM(4773) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4773)))) severity failure;
    assert RAM(4774) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4774)))) severity failure;
    assert RAM(4775) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4775)))) severity failure;
    assert RAM(4776) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4776)))) severity failure;
    assert RAM(4777) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4777)))) severity failure;
    assert RAM(4778) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4778)))) severity failure;
    assert RAM(4779) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4779)))) severity failure;
    assert RAM(4780) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4780)))) severity failure;
    assert RAM(4781) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4781)))) severity failure;
    assert RAM(4782) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4782)))) severity failure;
    assert RAM(4783) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4783)))) severity failure;
    assert RAM(4784) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4784)))) severity failure;
    assert RAM(4785) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4785)))) severity failure;
    assert RAM(4786) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4786)))) severity failure;
    assert RAM(4787) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4787)))) severity failure;
    assert RAM(4788) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4788)))) severity failure;
    assert RAM(4789) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4789)))) severity failure;
    assert RAM(4790) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4790)))) severity failure;
    assert RAM(4791) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4791)))) severity failure;
    assert RAM(4792) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4792)))) severity failure;
    assert RAM(4793) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4793)))) severity failure;
    assert RAM(4794) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4794)))) severity failure;
    assert RAM(4795) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4795)))) severity failure;
    assert RAM(4796) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4796)))) severity failure;
    assert RAM(4797) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4797)))) severity failure;
    assert RAM(4798) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4798)))) severity failure;
    assert RAM(4799) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4799)))) severity failure;
    assert RAM(4800) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4800)))) severity failure;
    assert RAM(4801) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4801)))) severity failure;
    assert RAM(4802) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4802)))) severity failure;
    assert RAM(4803) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4803)))) severity failure;
    assert RAM(4804) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4804)))) severity failure;
    assert RAM(4805) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4805)))) severity failure;
    assert RAM(4806) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4806)))) severity failure;
    assert RAM(4807) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4807)))) severity failure;
    assert RAM(4808) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4808)))) severity failure;
    assert RAM(4809) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4809)))) severity failure;
    assert RAM(4810) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4810)))) severity failure;
    assert RAM(4811) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4811)))) severity failure;
    assert RAM(4812) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4812)))) severity failure;
    assert RAM(4813) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4813)))) severity failure;
    assert RAM(4814) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4814)))) severity failure;
    assert RAM(4815) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4815)))) severity failure;
    assert RAM(4816) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4816)))) severity failure;
    assert RAM(4817) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4817)))) severity failure;
    assert RAM(4818) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4818)))) severity failure;
    assert RAM(4819) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4819)))) severity failure;
    assert RAM(4820) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4820)))) severity failure;
    assert RAM(4821) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4821)))) severity failure;
    assert RAM(4822) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4822)))) severity failure;
    assert RAM(4823) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4823)))) severity failure;
    assert RAM(4824) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4824)))) severity failure;
    assert RAM(4825) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4825)))) severity failure;
    assert RAM(4826) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4826)))) severity failure;
    assert RAM(4827) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4827)))) severity failure;
    assert RAM(4828) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4828)))) severity failure;
    assert RAM(4829) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4829)))) severity failure;
    assert RAM(4830) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4830)))) severity failure;
    assert RAM(4831) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4831)))) severity failure;
    assert RAM(4832) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4832)))) severity failure;
    assert RAM(4833) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4833)))) severity failure;
    assert RAM(4834) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4834)))) severity failure;
    assert RAM(4835) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4835)))) severity failure;
    assert RAM(4836) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4836)))) severity failure;
    assert RAM(4837) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4837)))) severity failure;
    assert RAM(4838) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4838)))) severity failure;
    assert RAM(4839) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4839)))) severity failure;
    assert RAM(4840) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4840)))) severity failure;
    assert RAM(4841) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4841)))) severity failure;
    assert RAM(4842) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4842)))) severity failure;
    assert RAM(4843) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4843)))) severity failure;
    assert RAM(4844) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4844)))) severity failure;
    assert RAM(4845) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4845)))) severity failure;
    assert RAM(4846) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4846)))) severity failure;
    assert RAM(4847) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4847)))) severity failure;
    assert RAM(4848) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4848)))) severity failure;
    assert RAM(4849) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4849)))) severity failure;
    assert RAM(4850) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4850)))) severity failure;
    assert RAM(4851) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4851)))) severity failure;
    assert RAM(4852) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4852)))) severity failure;
    assert RAM(4853) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4853)))) severity failure;
    assert RAM(4854) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4854)))) severity failure;
    assert RAM(4855) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4855)))) severity failure;
    assert RAM(4856) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4856)))) severity failure;
    assert RAM(4857) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4857)))) severity failure;
    assert RAM(4858) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4858)))) severity failure;
    assert RAM(4859) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4859)))) severity failure;
    assert RAM(4860) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4860)))) severity failure;
    assert RAM(4861) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4861)))) severity failure;
    assert RAM(4862) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4862)))) severity failure;
    assert RAM(4863) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4863)))) severity failure;
    assert RAM(4864) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4864)))) severity failure;
    assert RAM(4865) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4865)))) severity failure;
    assert RAM(4866) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4866)))) severity failure;
    assert RAM(4867) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4867)))) severity failure;
    assert RAM(4868) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4868)))) severity failure;
    assert RAM(4869) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4869)))) severity failure;
    assert RAM(4870) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4870)))) severity failure;
    assert RAM(4871) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4871)))) severity failure;
    assert RAM(4872) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4872)))) severity failure;
    assert RAM(4873) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4873)))) severity failure;
    assert RAM(4874) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4874)))) severity failure;
    assert RAM(4875) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4875)))) severity failure;
    assert RAM(4876) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4876)))) severity failure;
    assert RAM(4877) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4877)))) severity failure;
    assert RAM(4878) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4878)))) severity failure;
    assert RAM(4879) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4879)))) severity failure;
    assert RAM(4880) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4880)))) severity failure;
    assert RAM(4881) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4881)))) severity failure;
    assert RAM(4882) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4882)))) severity failure;
    assert RAM(4883) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4883)))) severity failure;
    assert RAM(4884) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4884)))) severity failure;
    assert RAM(4885) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4885)))) severity failure;
    assert RAM(4886) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4886)))) severity failure;
    assert RAM(4887) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4887)))) severity failure;
    assert RAM(4888) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4888)))) severity failure;
    assert RAM(4889) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4889)))) severity failure;
    assert RAM(4890) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4890)))) severity failure;
    assert RAM(4891) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4891)))) severity failure;
    assert RAM(4892) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4892)))) severity failure;
    assert RAM(4893) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4893)))) severity failure;
    assert RAM(4894) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4894)))) severity failure;
    assert RAM(4895) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4895)))) severity failure;
    assert RAM(4896) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4896)))) severity failure;
    assert RAM(4897) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4897)))) severity failure;
    assert RAM(4898) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4898)))) severity failure;
    assert RAM(4899) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4899)))) severity failure;
    assert RAM(4900) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4900)))) severity failure;
    assert RAM(4901) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4901)))) severity failure;
    assert RAM(4902) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4902)))) severity failure;
    assert RAM(4903) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4903)))) severity failure;
    assert RAM(4904) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4904)))) severity failure;
    assert RAM(4905) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4905)))) severity failure;
    assert RAM(4906) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4906)))) severity failure;
    assert RAM(4907) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4907)))) severity failure;
    assert RAM(4908) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4908)))) severity failure;
    assert RAM(4909) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4909)))) severity failure;
    assert RAM(4910) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4910)))) severity failure;
    assert RAM(4911) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4911)))) severity failure;
    assert RAM(4912) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4912)))) severity failure;
    assert RAM(4913) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4913)))) severity failure;
    assert RAM(4914) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4914)))) severity failure;
    assert RAM(4915) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4915)))) severity failure;
    assert RAM(4916) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4916)))) severity failure;
    assert RAM(4917) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4917)))) severity failure;
    assert RAM(4918) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4918)))) severity failure;
    assert RAM(4919) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4919)))) severity failure;
    assert RAM(4920) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4920)))) severity failure;
    assert RAM(4921) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4921)))) severity failure;
    assert RAM(4922) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4922)))) severity failure;
    assert RAM(4923) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4923)))) severity failure;
    assert RAM(4924) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4924)))) severity failure;
    assert RAM(4925) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4925)))) severity failure;
    assert RAM(4926) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4926)))) severity failure;
    assert RAM(4927) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4927)))) severity failure;
    assert RAM(4928) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4928)))) severity failure;
    assert RAM(4929) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4929)))) severity failure;
    assert RAM(4930) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4930)))) severity failure;
    assert RAM(4931) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4931)))) severity failure;
    assert RAM(4932) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4932)))) severity failure;
    assert RAM(4933) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4933)))) severity failure;
    assert RAM(4934) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4934)))) severity failure;
    assert RAM(4935) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4935)))) severity failure;
    assert RAM(4936) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4936)))) severity failure;
    assert RAM(4937) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4937)))) severity failure;
    assert RAM(4938) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4938)))) severity failure;
    assert RAM(4939) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4939)))) severity failure;
    assert RAM(4940) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4940)))) severity failure;
    assert RAM(4941) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4941)))) severity failure;
    assert RAM(4942) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4942)))) severity failure;
    assert RAM(4943) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4943)))) severity failure;
    assert RAM(4944) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4944)))) severity failure;
    assert RAM(4945) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4945)))) severity failure;
    assert RAM(4946) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4946)))) severity failure;
    assert RAM(4947) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4947)))) severity failure;
    assert RAM(4948) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4948)))) severity failure;
    assert RAM(4949) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4949)))) severity failure;
    assert RAM(4950) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4950)))) severity failure;
    assert RAM(4951) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4951)))) severity failure;
    assert RAM(4952) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4952)))) severity failure;
    assert RAM(4953) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4953)))) severity failure;
    assert RAM(4954) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4954)))) severity failure;
    assert RAM(4955) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4955)))) severity failure;
    assert RAM(4956) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4956)))) severity failure;
    assert RAM(4957) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4957)))) severity failure;
    assert RAM(4958) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4958)))) severity failure;
    assert RAM(4959) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4959)))) severity failure;
    assert RAM(4960) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4960)))) severity failure;
    assert RAM(4961) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4961)))) severity failure;
    assert RAM(4962) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4962)))) severity failure;
    assert RAM(4963) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4963)))) severity failure;
    assert RAM(4964) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4964)))) severity failure;
    assert RAM(4965) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4965)))) severity failure;
    assert RAM(4966) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(4966)))) severity failure;
    assert RAM(4967) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4967)))) severity failure;
    assert RAM(4968) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4968)))) severity failure;
    assert RAM(4969) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4969)))) severity failure;
    assert RAM(4970) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4970)))) severity failure;
    assert RAM(4971) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4971)))) severity failure;
    assert RAM(4972) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4972)))) severity failure;
    assert RAM(4973) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4973)))) severity failure;
    assert RAM(4974) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4974)))) severity failure;
    assert RAM(4975) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4975)))) severity failure;
    assert RAM(4976) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4976)))) severity failure;
    assert RAM(4977) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4977)))) severity failure;
    assert RAM(4978) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4978)))) severity failure;
    assert RAM(4979) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4979)))) severity failure;
    assert RAM(4980) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4980)))) severity failure;
    assert RAM(4981) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(4981)))) severity failure;
    assert RAM(4982) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4982)))) severity failure;
    assert RAM(4983) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4983)))) severity failure;
    assert RAM(4984) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(4984)))) severity failure;
    assert RAM(4985) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(4985)))) severity failure;
    assert RAM(4986) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4986)))) severity failure;
    assert RAM(4987) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4987)))) severity failure;
    assert RAM(4988) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4988)))) severity failure;
    assert RAM(4989) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(4989)))) severity failure;
    assert RAM(4990) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4990)))) severity failure;
    assert RAM(4991) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4991)))) severity failure;
    assert RAM(4992) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(4992)))) severity failure;
    assert RAM(4993) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4993)))) severity failure;
    assert RAM(4994) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4994)))) severity failure;
    assert RAM(4995) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4995)))) severity failure;
    assert RAM(4996) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4996)))) severity failure;
    assert RAM(4997) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(4997)))) severity failure;
    assert RAM(4998) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(4998)))) severity failure;
    assert RAM(4999) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(4999)))) severity failure;
    assert RAM(5000) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5000)))) severity failure;
    assert RAM(5001) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5001)))) severity failure;
    assert RAM(5002) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5002)))) severity failure;
    assert RAM(5003) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5003)))) severity failure;
    assert RAM(5004) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5004)))) severity failure;
    assert RAM(5005) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5005)))) severity failure;
    assert RAM(5006) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5006)))) severity failure;
    assert RAM(5007) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5007)))) severity failure;
    assert RAM(5008) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5008)))) severity failure;
    assert RAM(5009) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5009)))) severity failure;
    assert RAM(5010) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5010)))) severity failure;
    assert RAM(5011) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5011)))) severity failure;
    assert RAM(5012) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5012)))) severity failure;
    assert RAM(5013) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5013)))) severity failure;
    assert RAM(5014) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5014)))) severity failure;
    assert RAM(5015) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5015)))) severity failure;
    assert RAM(5016) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5016)))) severity failure;
    assert RAM(5017) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5017)))) severity failure;
    assert RAM(5018) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5018)))) severity failure;
    assert RAM(5019) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5019)))) severity failure;
    assert RAM(5020) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5020)))) severity failure;
    assert RAM(5021) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5021)))) severity failure;
    assert RAM(5022) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5022)))) severity failure;
    assert RAM(5023) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5023)))) severity failure;
    assert RAM(5024) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5024)))) severity failure;
    assert RAM(5025) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5025)))) severity failure;
    assert RAM(5026) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5026)))) severity failure;
    assert RAM(5027) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5027)))) severity failure;
    assert RAM(5028) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5028)))) severity failure;
    assert RAM(5029) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5029)))) severity failure;
    assert RAM(5030) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5030)))) severity failure;
    assert RAM(5031) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5031)))) severity failure;
    assert RAM(5032) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5032)))) severity failure;
    assert RAM(5033) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5033)))) severity failure;
    assert RAM(5034) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5034)))) severity failure;
    assert RAM(5035) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5035)))) severity failure;
    assert RAM(5036) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5036)))) severity failure;
    assert RAM(5037) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5037)))) severity failure;
    assert RAM(5038) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5038)))) severity failure;
    assert RAM(5039) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5039)))) severity failure;
    assert RAM(5040) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5040)))) severity failure;
    assert RAM(5041) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5041)))) severity failure;
    assert RAM(5042) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5042)))) severity failure;
    assert RAM(5043) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5043)))) severity failure;
    assert RAM(5044) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5044)))) severity failure;
    assert RAM(5045) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5045)))) severity failure;
    assert RAM(5046) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5046)))) severity failure;
    assert RAM(5047) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5047)))) severity failure;
    assert RAM(5048) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5048)))) severity failure;
    assert RAM(5049) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5049)))) severity failure;
    assert RAM(5050) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5050)))) severity failure;
    assert RAM(5051) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5051)))) severity failure;
    assert RAM(5052) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5052)))) severity failure;
    assert RAM(5053) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5053)))) severity failure;
    assert RAM(5054) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5054)))) severity failure;
    assert RAM(5055) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5055)))) severity failure;
    assert RAM(5056) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5056)))) severity failure;
    assert RAM(5057) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5057)))) severity failure;
    assert RAM(5058) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5058)))) severity failure;
    assert RAM(5059) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5059)))) severity failure;
    assert RAM(5060) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5060)))) severity failure;
    assert RAM(5061) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5061)))) severity failure;
    assert RAM(5062) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5062)))) severity failure;
    assert RAM(5063) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5063)))) severity failure;
    assert RAM(5064) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5064)))) severity failure;
    assert RAM(5065) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5065)))) severity failure;
    assert RAM(5066) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5066)))) severity failure;
    assert RAM(5067) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5067)))) severity failure;
    assert RAM(5068) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5068)))) severity failure;
    assert RAM(5069) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5069)))) severity failure;
    assert RAM(5070) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5070)))) severity failure;
    assert RAM(5071) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5071)))) severity failure;
    assert RAM(5072) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5072)))) severity failure;
    assert RAM(5073) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5073)))) severity failure;
    assert RAM(5074) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5074)))) severity failure;
    assert RAM(5075) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5075)))) severity failure;
    assert RAM(5076) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5076)))) severity failure;
    assert RAM(5077) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5077)))) severity failure;
    assert RAM(5078) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5078)))) severity failure;
    assert RAM(5079) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5079)))) severity failure;
    assert RAM(5080) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5080)))) severity failure;
    assert RAM(5081) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5081)))) severity failure;
    assert RAM(5082) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5082)))) severity failure;
    assert RAM(5083) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5083)))) severity failure;
    assert RAM(5084) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5084)))) severity failure;
    assert RAM(5085) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5085)))) severity failure;
    assert RAM(5086) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5086)))) severity failure;
    assert RAM(5087) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5087)))) severity failure;
    assert RAM(5088) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5088)))) severity failure;
    assert RAM(5089) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5089)))) severity failure;
    assert RAM(5090) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5090)))) severity failure;
    assert RAM(5091) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5091)))) severity failure;
    assert RAM(5092) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5092)))) severity failure;
    assert RAM(5093) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5093)))) severity failure;
    assert RAM(5094) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5094)))) severity failure;
    assert RAM(5095) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5095)))) severity failure;
    assert RAM(5096) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5096)))) severity failure;
    assert RAM(5097) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5097)))) severity failure;
    assert RAM(5098) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5098)))) severity failure;
    assert RAM(5099) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5099)))) severity failure;
    assert RAM(5100) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5100)))) severity failure;
    assert RAM(5101) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5101)))) severity failure;
    assert RAM(5102) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5102)))) severity failure;
    assert RAM(5103) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5103)))) severity failure;
    assert RAM(5104) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5104)))) severity failure;
    assert RAM(5105) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5105)))) severity failure;
    assert RAM(5106) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5106)))) severity failure;
    assert RAM(5107) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5107)))) severity failure;
    assert RAM(5108) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5108)))) severity failure;
    assert RAM(5109) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5109)))) severity failure;
    assert RAM(5110) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5110)))) severity failure;
    assert RAM(5111) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5111)))) severity failure;
    assert RAM(5112) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5112)))) severity failure;
    assert RAM(5113) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5113)))) severity failure;
    assert RAM(5114) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5114)))) severity failure;
    assert RAM(5115) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5115)))) severity failure;
    assert RAM(5116) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5116)))) severity failure;
    assert RAM(5117) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5117)))) severity failure;
    assert RAM(5118) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5118)))) severity failure;
    assert RAM(5119) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5119)))) severity failure;
    assert RAM(5120) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5120)))) severity failure;
    assert RAM(5121) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5121)))) severity failure;
    assert RAM(5122) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5122)))) severity failure;
    assert RAM(5123) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5123)))) severity failure;
    assert RAM(5124) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5124)))) severity failure;
    assert RAM(5125) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5125)))) severity failure;
    assert RAM(5126) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5126)))) severity failure;
    assert RAM(5127) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5127)))) severity failure;
    assert RAM(5128) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5128)))) severity failure;
    assert RAM(5129) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5129)))) severity failure;
    assert RAM(5130) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5130)))) severity failure;
    assert RAM(5131) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5131)))) severity failure;
    assert RAM(5132) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5132)))) severity failure;
    assert RAM(5133) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5133)))) severity failure;
    assert RAM(5134) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5134)))) severity failure;
    assert RAM(5135) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5135)))) severity failure;
    assert RAM(5136) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5136)))) severity failure;
    assert RAM(5137) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5137)))) severity failure;
    assert RAM(5138) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5138)))) severity failure;
    assert RAM(5139) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5139)))) severity failure;
    assert RAM(5140) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5140)))) severity failure;
    assert RAM(5141) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5141)))) severity failure;
    assert RAM(5142) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5142)))) severity failure;
    assert RAM(5143) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5143)))) severity failure;
    assert RAM(5144) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5144)))) severity failure;
    assert RAM(5145) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5145)))) severity failure;
    assert RAM(5146) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5146)))) severity failure;
    assert RAM(5147) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5147)))) severity failure;
    assert RAM(5148) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5148)))) severity failure;
    assert RAM(5149) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5149)))) severity failure;
    assert RAM(5150) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5150)))) severity failure;
    assert RAM(5151) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5151)))) severity failure;
    assert RAM(5152) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5152)))) severity failure;
    assert RAM(5153) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5153)))) severity failure;
    assert RAM(5154) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5154)))) severity failure;
    assert RAM(5155) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5155)))) severity failure;
    assert RAM(5156) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5156)))) severity failure;
    assert RAM(5157) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5157)))) severity failure;
    assert RAM(5158) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5158)))) severity failure;
    assert RAM(5159) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5159)))) severity failure;
    assert RAM(5160) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5160)))) severity failure;
    assert RAM(5161) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5161)))) severity failure;
    assert RAM(5162) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5162)))) severity failure;
    assert RAM(5163) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5163)))) severity failure;
    assert RAM(5164) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5164)))) severity failure;
    assert RAM(5165) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5165)))) severity failure;
    assert RAM(5166) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5166)))) severity failure;
    assert RAM(5167) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5167)))) severity failure;
    assert RAM(5168) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5168)))) severity failure;
    assert RAM(5169) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5169)))) severity failure;
    assert RAM(5170) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5170)))) severity failure;
    assert RAM(5171) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5171)))) severity failure;
    assert RAM(5172) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5172)))) severity failure;
    assert RAM(5173) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5173)))) severity failure;
    assert RAM(5174) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5174)))) severity failure;
    assert RAM(5175) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5175)))) severity failure;
    assert RAM(5176) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5176)))) severity failure;
    assert RAM(5177) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5177)))) severity failure;
    assert RAM(5178) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5178)))) severity failure;
    assert RAM(5179) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5179)))) severity failure;
    assert RAM(5180) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5180)))) severity failure;
    assert RAM(5181) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5181)))) severity failure;
    assert RAM(5182) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5182)))) severity failure;
    assert RAM(5183) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5183)))) severity failure;
    assert RAM(5184) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5184)))) severity failure;
    assert RAM(5185) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5185)))) severity failure;
    assert RAM(5186) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5186)))) severity failure;
    assert RAM(5187) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5187)))) severity failure;
    assert RAM(5188) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5188)))) severity failure;
    assert RAM(5189) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5189)))) severity failure;
    assert RAM(5190) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5190)))) severity failure;
    assert RAM(5191) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5191)))) severity failure;
    assert RAM(5192) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5192)))) severity failure;
    assert RAM(5193) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5193)))) severity failure;
    assert RAM(5194) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5194)))) severity failure;
    assert RAM(5195) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5195)))) severity failure;
    assert RAM(5196) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5196)))) severity failure;
    assert RAM(5197) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5197)))) severity failure;
    assert RAM(5198) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5198)))) severity failure;
    assert RAM(5199) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5199)))) severity failure;
    assert RAM(5200) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5200)))) severity failure;
    assert RAM(5201) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5201)))) severity failure;
    assert RAM(5202) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5202)))) severity failure;
    assert RAM(5203) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5203)))) severity failure;
    assert RAM(5204) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5204)))) severity failure;
    assert RAM(5205) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5205)))) severity failure;
    assert RAM(5206) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5206)))) severity failure;
    assert RAM(5207) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5207)))) severity failure;
    assert RAM(5208) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5208)))) severity failure;
    assert RAM(5209) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5209)))) severity failure;
    assert RAM(5210) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5210)))) severity failure;
    assert RAM(5211) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5211)))) severity failure;
    assert RAM(5212) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5212)))) severity failure;
    assert RAM(5213) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5213)))) severity failure;
    assert RAM(5214) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5214)))) severity failure;
    assert RAM(5215) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5215)))) severity failure;
    assert RAM(5216) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5216)))) severity failure;
    assert RAM(5217) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5217)))) severity failure;
    assert RAM(5218) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5218)))) severity failure;
    assert RAM(5219) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5219)))) severity failure;
    assert RAM(5220) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5220)))) severity failure;
    assert RAM(5221) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5221)))) severity failure;
    assert RAM(5222) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5222)))) severity failure;
    assert RAM(5223) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5223)))) severity failure;
    assert RAM(5224) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5224)))) severity failure;
    assert RAM(5225) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5225)))) severity failure;
    assert RAM(5226) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5226)))) severity failure;
    assert RAM(5227) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5227)))) severity failure;
    assert RAM(5228) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5228)))) severity failure;
    assert RAM(5229) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5229)))) severity failure;
    assert RAM(5230) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5230)))) severity failure;
    assert RAM(5231) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5231)))) severity failure;
    assert RAM(5232) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5232)))) severity failure;
    assert RAM(5233) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5233)))) severity failure;
    assert RAM(5234) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5234)))) severity failure;
    assert RAM(5235) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5235)))) severity failure;
    assert RAM(5236) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5236)))) severity failure;
    assert RAM(5237) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5237)))) severity failure;
    assert RAM(5238) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5238)))) severity failure;
    assert RAM(5239) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5239)))) severity failure;
    assert RAM(5240) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5240)))) severity failure;
    assert RAM(5241) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5241)))) severity failure;
    assert RAM(5242) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5242)))) severity failure;
    assert RAM(5243) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5243)))) severity failure;
    assert RAM(5244) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5244)))) severity failure;
    assert RAM(5245) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5245)))) severity failure;
    assert RAM(5246) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5246)))) severity failure;
    assert RAM(5247) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5247)))) severity failure;
    assert RAM(5248) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5248)))) severity failure;
    assert RAM(5249) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5249)))) severity failure;
    assert RAM(5250) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5250)))) severity failure;
    assert RAM(5251) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5251)))) severity failure;
    assert RAM(5252) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5252)))) severity failure;
    assert RAM(5253) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5253)))) severity failure;
    assert RAM(5254) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5254)))) severity failure;
    assert RAM(5255) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5255)))) severity failure;
    assert RAM(5256) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5256)))) severity failure;
    assert RAM(5257) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5257)))) severity failure;
    assert RAM(5258) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5258)))) severity failure;
    assert RAM(5259) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5259)))) severity failure;
    assert RAM(5260) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5260)))) severity failure;
    assert RAM(5261) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5261)))) severity failure;
    assert RAM(5262) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5262)))) severity failure;
    assert RAM(5263) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5263)))) severity failure;
    assert RAM(5264) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5264)))) severity failure;
    assert RAM(5265) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5265)))) severity failure;
    assert RAM(5266) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5266)))) severity failure;
    assert RAM(5267) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5267)))) severity failure;
    assert RAM(5268) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5268)))) severity failure;
    assert RAM(5269) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5269)))) severity failure;
    assert RAM(5270) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5270)))) severity failure;
    assert RAM(5271) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5271)))) severity failure;
    assert RAM(5272) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5272)))) severity failure;
    assert RAM(5273) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5273)))) severity failure;
    assert RAM(5274) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5274)))) severity failure;
    assert RAM(5275) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5275)))) severity failure;
    assert RAM(5276) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5276)))) severity failure;
    assert RAM(5277) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5277)))) severity failure;
    assert RAM(5278) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5278)))) severity failure;
    assert RAM(5279) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5279)))) severity failure;
    assert RAM(5280) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5280)))) severity failure;
    assert RAM(5281) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5281)))) severity failure;
    assert RAM(5282) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5282)))) severity failure;
    assert RAM(5283) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5283)))) severity failure;
    assert RAM(5284) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5284)))) severity failure;
    assert RAM(5285) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5285)))) severity failure;
    assert RAM(5286) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5286)))) severity failure;
    assert RAM(5287) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5287)))) severity failure;
    assert RAM(5288) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5288)))) severity failure;
    assert RAM(5289) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5289)))) severity failure;
    assert RAM(5290) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5290)))) severity failure;
    assert RAM(5291) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5291)))) severity failure;
    assert RAM(5292) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5292)))) severity failure;
    assert RAM(5293) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5293)))) severity failure;
    assert RAM(5294) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5294)))) severity failure;
    assert RAM(5295) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5295)))) severity failure;
    assert RAM(5296) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5296)))) severity failure;
    assert RAM(5297) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5297)))) severity failure;
    assert RAM(5298) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5298)))) severity failure;
    assert RAM(5299) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5299)))) severity failure;
    assert RAM(5300) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5300)))) severity failure;
    assert RAM(5301) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5301)))) severity failure;
    assert RAM(5302) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5302)))) severity failure;
    assert RAM(5303) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5303)))) severity failure;
    assert RAM(5304) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5304)))) severity failure;
    assert RAM(5305) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5305)))) severity failure;
    assert RAM(5306) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5306)))) severity failure;
    assert RAM(5307) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5307)))) severity failure;
    assert RAM(5308) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5308)))) severity failure;
    assert RAM(5309) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5309)))) severity failure;
    assert RAM(5310) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5310)))) severity failure;
    assert RAM(5311) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5311)))) severity failure;
    assert RAM(5312) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5312)))) severity failure;
    assert RAM(5313) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5313)))) severity failure;
    assert RAM(5314) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5314)))) severity failure;
    assert RAM(5315) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5315)))) severity failure;
    assert RAM(5316) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5316)))) severity failure;
    assert RAM(5317) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5317)))) severity failure;
    assert RAM(5318) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5318)))) severity failure;
    assert RAM(5319) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5319)))) severity failure;
    assert RAM(5320) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5320)))) severity failure;
    assert RAM(5321) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5321)))) severity failure;
    assert RAM(5322) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5322)))) severity failure;
    assert RAM(5323) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5323)))) severity failure;
    assert RAM(5324) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5324)))) severity failure;
    assert RAM(5325) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5325)))) severity failure;
    assert RAM(5326) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5326)))) severity failure;
    assert RAM(5327) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5327)))) severity failure;
    assert RAM(5328) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5328)))) severity failure;
    assert RAM(5329) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5329)))) severity failure;
    assert RAM(5330) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5330)))) severity failure;
    assert RAM(5331) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5331)))) severity failure;
    assert RAM(5332) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5332)))) severity failure;
    assert RAM(5333) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5333)))) severity failure;
    assert RAM(5334) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5334)))) severity failure;
    assert RAM(5335) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5335)))) severity failure;
    assert RAM(5336) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5336)))) severity failure;
    assert RAM(5337) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5337)))) severity failure;
    assert RAM(5338) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5338)))) severity failure;
    assert RAM(5339) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5339)))) severity failure;
    assert RAM(5340) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5340)))) severity failure;
    assert RAM(5341) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5341)))) severity failure;
    assert RAM(5342) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5342)))) severity failure;
    assert RAM(5343) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5343)))) severity failure;
    assert RAM(5344) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5344)))) severity failure;
    assert RAM(5345) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5345)))) severity failure;
    assert RAM(5346) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5346)))) severity failure;
    assert RAM(5347) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5347)))) severity failure;
    assert RAM(5348) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5348)))) severity failure;
    assert RAM(5349) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5349)))) severity failure;
    assert RAM(5350) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5350)))) severity failure;
    assert RAM(5351) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5351)))) severity failure;
    assert RAM(5352) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5352)))) severity failure;
    assert RAM(5353) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5353)))) severity failure;
    assert RAM(5354) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5354)))) severity failure;
    assert RAM(5355) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5355)))) severity failure;
    assert RAM(5356) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5356)))) severity failure;
    assert RAM(5357) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5357)))) severity failure;
    assert RAM(5358) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5358)))) severity failure;
    assert RAM(5359) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5359)))) severity failure;
    assert RAM(5360) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5360)))) severity failure;
    assert RAM(5361) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5361)))) severity failure;
    assert RAM(5362) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5362)))) severity failure;
    assert RAM(5363) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5363)))) severity failure;
    assert RAM(5364) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5364)))) severity failure;
    assert RAM(5365) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5365)))) severity failure;
    assert RAM(5366) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5366)))) severity failure;
    assert RAM(5367) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5367)))) severity failure;
    assert RAM(5368) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5368)))) severity failure;
    assert RAM(5369) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5369)))) severity failure;
    assert RAM(5370) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5370)))) severity failure;
    assert RAM(5371) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5371)))) severity failure;
    assert RAM(5372) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5372)))) severity failure;
    assert RAM(5373) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5373)))) severity failure;
    assert RAM(5374) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5374)))) severity failure;
    assert RAM(5375) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5375)))) severity failure;
    assert RAM(5376) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5376)))) severity failure;
    assert RAM(5377) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5377)))) severity failure;
    assert RAM(5378) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5378)))) severity failure;
    assert RAM(5379) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5379)))) severity failure;
    assert RAM(5380) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5380)))) severity failure;
    assert RAM(5381) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5381)))) severity failure;
    assert RAM(5382) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5382)))) severity failure;
    assert RAM(5383) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5383)))) severity failure;
    assert RAM(5384) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5384)))) severity failure;
    assert RAM(5385) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5385)))) severity failure;
    assert RAM(5386) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5386)))) severity failure;
    assert RAM(5387) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5387)))) severity failure;
    assert RAM(5388) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5388)))) severity failure;
    assert RAM(5389) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5389)))) severity failure;
    assert RAM(5390) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5390)))) severity failure;
    assert RAM(5391) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5391)))) severity failure;
    assert RAM(5392) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5392)))) severity failure;
    assert RAM(5393) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5393)))) severity failure;
    assert RAM(5394) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5394)))) severity failure;
    assert RAM(5395) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5395)))) severity failure;
    assert RAM(5396) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5396)))) severity failure;
    assert RAM(5397) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5397)))) severity failure;
    assert RAM(5398) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5398)))) severity failure;
    assert RAM(5399) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5399)))) severity failure;
    assert RAM(5400) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5400)))) severity failure;
    assert RAM(5401) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5401)))) severity failure;
    assert RAM(5402) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5402)))) severity failure;
    assert RAM(5403) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5403)))) severity failure;
    assert RAM(5404) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5404)))) severity failure;
    assert RAM(5405) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5405)))) severity failure;
    assert RAM(5406) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5406)))) severity failure;
    assert RAM(5407) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5407)))) severity failure;
    assert RAM(5408) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5408)))) severity failure;
    assert RAM(5409) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5409)))) severity failure;
    assert RAM(5410) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5410)))) severity failure;
    assert RAM(5411) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5411)))) severity failure;
    assert RAM(5412) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5412)))) severity failure;
    assert RAM(5413) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5413)))) severity failure;
    assert RAM(5414) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5414)))) severity failure;
    assert RAM(5415) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5415)))) severity failure;
    assert RAM(5416) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5416)))) severity failure;
    assert RAM(5417) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5417)))) severity failure;
    assert RAM(5418) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5418)))) severity failure;
    assert RAM(5419) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5419)))) severity failure;
    assert RAM(5420) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5420)))) severity failure;
    assert RAM(5421) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5421)))) severity failure;
    assert RAM(5422) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5422)))) severity failure;
    assert RAM(5423) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5423)))) severity failure;
    assert RAM(5424) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5424)))) severity failure;
    assert RAM(5425) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5425)))) severity failure;
    assert RAM(5426) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5426)))) severity failure;
    assert RAM(5427) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5427)))) severity failure;
    assert RAM(5428) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5428)))) severity failure;
    assert RAM(5429) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5429)))) severity failure;
    assert RAM(5430) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5430)))) severity failure;
    assert RAM(5431) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5431)))) severity failure;
    assert RAM(5432) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5432)))) severity failure;
    assert RAM(5433) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5433)))) severity failure;
    assert RAM(5434) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5434)))) severity failure;
    assert RAM(5435) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5435)))) severity failure;
    assert RAM(5436) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5436)))) severity failure;
    assert RAM(5437) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5437)))) severity failure;
    assert RAM(5438) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5438)))) severity failure;
    assert RAM(5439) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5439)))) severity failure;
    assert RAM(5440) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5440)))) severity failure;
    assert RAM(5441) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5441)))) severity failure;
    assert RAM(5442) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5442)))) severity failure;
    assert RAM(5443) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5443)))) severity failure;
    assert RAM(5444) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5444)))) severity failure;
    assert RAM(5445) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5445)))) severity failure;
    assert RAM(5446) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5446)))) severity failure;
    assert RAM(5447) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5447)))) severity failure;
    assert RAM(5448) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5448)))) severity failure;
    assert RAM(5449) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5449)))) severity failure;
    assert RAM(5450) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5450)))) severity failure;
    assert RAM(5451) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5451)))) severity failure;
    assert RAM(5452) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5452)))) severity failure;
    assert RAM(5453) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5453)))) severity failure;
    assert RAM(5454) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5454)))) severity failure;
    assert RAM(5455) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5455)))) severity failure;
    assert RAM(5456) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5456)))) severity failure;
    assert RAM(5457) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5457)))) severity failure;
    assert RAM(5458) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5458)))) severity failure;
    assert RAM(5459) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5459)))) severity failure;
    assert RAM(5460) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5460)))) severity failure;
    assert RAM(5461) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5461)))) severity failure;
    assert RAM(5462) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5462)))) severity failure;
    assert RAM(5463) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5463)))) severity failure;
    assert RAM(5464) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5464)))) severity failure;
    assert RAM(5465) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5465)))) severity failure;
    assert RAM(5466) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5466)))) severity failure;
    assert RAM(5467) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5467)))) severity failure;
    assert RAM(5468) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5468)))) severity failure;
    assert RAM(5469) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5469)))) severity failure;
    assert RAM(5470) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5470)))) severity failure;
    assert RAM(5471) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5471)))) severity failure;
    assert RAM(5472) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5472)))) severity failure;
    assert RAM(5473) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5473)))) severity failure;
    assert RAM(5474) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5474)))) severity failure;
    assert RAM(5475) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5475)))) severity failure;
    assert RAM(5476) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5476)))) severity failure;
    assert RAM(5477) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5477)))) severity failure;
    assert RAM(5478) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5478)))) severity failure;
    assert RAM(5479) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5479)))) severity failure;
    assert RAM(5480) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5480)))) severity failure;
    assert RAM(5481) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5481)))) severity failure;
    assert RAM(5482) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5482)))) severity failure;
    assert RAM(5483) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5483)))) severity failure;
    assert RAM(5484) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5484)))) severity failure;
    assert RAM(5485) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5485)))) severity failure;
    assert RAM(5486) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5486)))) severity failure;
    assert RAM(5487) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5487)))) severity failure;
    assert RAM(5488) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5488)))) severity failure;
    assert RAM(5489) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5489)))) severity failure;
    assert RAM(5490) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5490)))) severity failure;
    assert RAM(5491) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5491)))) severity failure;
    assert RAM(5492) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5492)))) severity failure;
    assert RAM(5493) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5493)))) severity failure;
    assert RAM(5494) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5494)))) severity failure;
    assert RAM(5495) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5495)))) severity failure;
    assert RAM(5496) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5496)))) severity failure;
    assert RAM(5497) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5497)))) severity failure;
    assert RAM(5498) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5498)))) severity failure;
    assert RAM(5499) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5499)))) severity failure;
    assert RAM(5500) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5500)))) severity failure;
    assert RAM(5501) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5501)))) severity failure;
    assert RAM(5502) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5502)))) severity failure;
    assert RAM(5503) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5503)))) severity failure;
    assert RAM(5504) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5504)))) severity failure;
    assert RAM(5505) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5505)))) severity failure;
    assert RAM(5506) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5506)))) severity failure;
    assert RAM(5507) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5507)))) severity failure;
    assert RAM(5508) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5508)))) severity failure;
    assert RAM(5509) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5509)))) severity failure;
    assert RAM(5510) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5510)))) severity failure;
    assert RAM(5511) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5511)))) severity failure;
    assert RAM(5512) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5512)))) severity failure;
    assert RAM(5513) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5513)))) severity failure;
    assert RAM(5514) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5514)))) severity failure;
    assert RAM(5515) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5515)))) severity failure;
    assert RAM(5516) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5516)))) severity failure;
    assert RAM(5517) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5517)))) severity failure;
    assert RAM(5518) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5518)))) severity failure;
    assert RAM(5519) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5519)))) severity failure;
    assert RAM(5520) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5520)))) severity failure;
    assert RAM(5521) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5521)))) severity failure;
    assert RAM(5522) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5522)))) severity failure;
    assert RAM(5523) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5523)))) severity failure;
    assert RAM(5524) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5524)))) severity failure;
    assert RAM(5525) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5525)))) severity failure;
    assert RAM(5526) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5526)))) severity failure;
    assert RAM(5527) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5527)))) severity failure;
    assert RAM(5528) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5528)))) severity failure;
    assert RAM(5529) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5529)))) severity failure;
    assert RAM(5530) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5530)))) severity failure;
    assert RAM(5531) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5531)))) severity failure;
    assert RAM(5532) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5532)))) severity failure;
    assert RAM(5533) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5533)))) severity failure;
    assert RAM(5534) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5534)))) severity failure;
    assert RAM(5535) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5535)))) severity failure;
    assert RAM(5536) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5536)))) severity failure;
    assert RAM(5537) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5537)))) severity failure;
    assert RAM(5538) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5538)))) severity failure;
    assert RAM(5539) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5539)))) severity failure;
    assert RAM(5540) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5540)))) severity failure;
    assert RAM(5541) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5541)))) severity failure;
    assert RAM(5542) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5542)))) severity failure;
    assert RAM(5543) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5543)))) severity failure;
    assert RAM(5544) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5544)))) severity failure;
    assert RAM(5545) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5545)))) severity failure;
    assert RAM(5546) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5546)))) severity failure;
    assert RAM(5547) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5547)))) severity failure;
    assert RAM(5548) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5548)))) severity failure;
    assert RAM(5549) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5549)))) severity failure;
    assert RAM(5550) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5550)))) severity failure;
    assert RAM(5551) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5551)))) severity failure;
    assert RAM(5552) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5552)))) severity failure;
    assert RAM(5553) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5553)))) severity failure;
    assert RAM(5554) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5554)))) severity failure;
    assert RAM(5555) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5555)))) severity failure;
    assert RAM(5556) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5556)))) severity failure;
    assert RAM(5557) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5557)))) severity failure;
    assert RAM(5558) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5558)))) severity failure;
    assert RAM(5559) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5559)))) severity failure;
    assert RAM(5560) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5560)))) severity failure;
    assert RAM(5561) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5561)))) severity failure;
    assert RAM(5562) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5562)))) severity failure;
    assert RAM(5563) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5563)))) severity failure;
    assert RAM(5564) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5564)))) severity failure;
    assert RAM(5565) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5565)))) severity failure;
    assert RAM(5566) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5566)))) severity failure;
    assert RAM(5567) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5567)))) severity failure;
    assert RAM(5568) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5568)))) severity failure;
    assert RAM(5569) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5569)))) severity failure;
    assert RAM(5570) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5570)))) severity failure;
    assert RAM(5571) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5571)))) severity failure;
    assert RAM(5572) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5572)))) severity failure;
    assert RAM(5573) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5573)))) severity failure;
    assert RAM(5574) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5574)))) severity failure;
    assert RAM(5575) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5575)))) severity failure;
    assert RAM(5576) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5576)))) severity failure;
    assert RAM(5577) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5577)))) severity failure;
    assert RAM(5578) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5578)))) severity failure;
    assert RAM(5579) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5579)))) severity failure;
    assert RAM(5580) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5580)))) severity failure;
    assert RAM(5581) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5581)))) severity failure;
    assert RAM(5582) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5582)))) severity failure;
    assert RAM(5583) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5583)))) severity failure;
    assert RAM(5584) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5584)))) severity failure;
    assert RAM(5585) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5585)))) severity failure;
    assert RAM(5586) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5586)))) severity failure;
    assert RAM(5587) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5587)))) severity failure;
    assert RAM(5588) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5588)))) severity failure;
    assert RAM(5589) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5589)))) severity failure;
    assert RAM(5590) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5590)))) severity failure;
    assert RAM(5591) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5591)))) severity failure;
    assert RAM(5592) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5592)))) severity failure;
    assert RAM(5593) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5593)))) severity failure;
    assert RAM(5594) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5594)))) severity failure;
    assert RAM(5595) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5595)))) severity failure;
    assert RAM(5596) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5596)))) severity failure;
    assert RAM(5597) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5597)))) severity failure;
    assert RAM(5598) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5598)))) severity failure;
    assert RAM(5599) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5599)))) severity failure;
    assert RAM(5600) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5600)))) severity failure;
    assert RAM(5601) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5601)))) severity failure;
    assert RAM(5602) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5602)))) severity failure;
    assert RAM(5603) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5603)))) severity failure;
    assert RAM(5604) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5604)))) severity failure;
    assert RAM(5605) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5605)))) severity failure;
    assert RAM(5606) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5606)))) severity failure;
    assert RAM(5607) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5607)))) severity failure;
    assert RAM(5608) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5608)))) severity failure;
    assert RAM(5609) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5609)))) severity failure;
    assert RAM(5610) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5610)))) severity failure;
    assert RAM(5611) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5611)))) severity failure;
    assert RAM(5612) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5612)))) severity failure;
    assert RAM(5613) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5613)))) severity failure;
    assert RAM(5614) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5614)))) severity failure;
    assert RAM(5615) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5615)))) severity failure;
    assert RAM(5616) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5616)))) severity failure;
    assert RAM(5617) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5617)))) severity failure;
    assert RAM(5618) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5618)))) severity failure;
    assert RAM(5619) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5619)))) severity failure;
    assert RAM(5620) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5620)))) severity failure;
    assert RAM(5621) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5621)))) severity failure;
    assert RAM(5622) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5622)))) severity failure;
    assert RAM(5623) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5623)))) severity failure;
    assert RAM(5624) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5624)))) severity failure;
    assert RAM(5625) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5625)))) severity failure;
    assert RAM(5626) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5626)))) severity failure;
    assert RAM(5627) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5627)))) severity failure;
    assert RAM(5628) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5628)))) severity failure;
    assert RAM(5629) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5629)))) severity failure;
    assert RAM(5630) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5630)))) severity failure;
    assert RAM(5631) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5631)))) severity failure;
    assert RAM(5632) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5632)))) severity failure;
    assert RAM(5633) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5633)))) severity failure;
    assert RAM(5634) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5634)))) severity failure;
    assert RAM(5635) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5635)))) severity failure;
    assert RAM(5636) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5636)))) severity failure;
    assert RAM(5637) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5637)))) severity failure;
    assert RAM(5638) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5638)))) severity failure;
    assert RAM(5639) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5639)))) severity failure;
    assert RAM(5640) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5640)))) severity failure;
    assert RAM(5641) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5641)))) severity failure;
    assert RAM(5642) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5642)))) severity failure;
    assert RAM(5643) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5643)))) severity failure;
    assert RAM(5644) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5644)))) severity failure;
    assert RAM(5645) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5645)))) severity failure;
    assert RAM(5646) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5646)))) severity failure;
    assert RAM(5647) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5647)))) severity failure;
    assert RAM(5648) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5648)))) severity failure;
    assert RAM(5649) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5649)))) severity failure;
    assert RAM(5650) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5650)))) severity failure;
    assert RAM(5651) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5651)))) severity failure;
    assert RAM(5652) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5652)))) severity failure;
    assert RAM(5653) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5653)))) severity failure;
    assert RAM(5654) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5654)))) severity failure;
    assert RAM(5655) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5655)))) severity failure;
    assert RAM(5656) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5656)))) severity failure;
    assert RAM(5657) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5657)))) severity failure;
    assert RAM(5658) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5658)))) severity failure;
    assert RAM(5659) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5659)))) severity failure;
    assert RAM(5660) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5660)))) severity failure;
    assert RAM(5661) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5661)))) severity failure;
    assert RAM(5662) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5662)))) severity failure;
    assert RAM(5663) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5663)))) severity failure;
    assert RAM(5664) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5664)))) severity failure;
    assert RAM(5665) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5665)))) severity failure;
    assert RAM(5666) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5666)))) severity failure;
    assert RAM(5667) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5667)))) severity failure;
    assert RAM(5668) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5668)))) severity failure;
    assert RAM(5669) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5669)))) severity failure;
    assert RAM(5670) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5670)))) severity failure;
    assert RAM(5671) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5671)))) severity failure;
    assert RAM(5672) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5672)))) severity failure;
    assert RAM(5673) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5673)))) severity failure;
    assert RAM(5674) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5674)))) severity failure;
    assert RAM(5675) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5675)))) severity failure;
    assert RAM(5676) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5676)))) severity failure;
    assert RAM(5677) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5677)))) severity failure;
    assert RAM(5678) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5678)))) severity failure;
    assert RAM(5679) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5679)))) severity failure;
    assert RAM(5680) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5680)))) severity failure;
    assert RAM(5681) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5681)))) severity failure;
    assert RAM(5682) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5682)))) severity failure;
    assert RAM(5683) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5683)))) severity failure;
    assert RAM(5684) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5684)))) severity failure;
    assert RAM(5685) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5685)))) severity failure;
    assert RAM(5686) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5686)))) severity failure;
    assert RAM(5687) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5687)))) severity failure;
    assert RAM(5688) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5688)))) severity failure;
    assert RAM(5689) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5689)))) severity failure;
    assert RAM(5690) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5690)))) severity failure;
    assert RAM(5691) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5691)))) severity failure;
    assert RAM(5692) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5692)))) severity failure;
    assert RAM(5693) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5693)))) severity failure;
    assert RAM(5694) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5694)))) severity failure;
    assert RAM(5695) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5695)))) severity failure;
    assert RAM(5696) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5696)))) severity failure;
    assert RAM(5697) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5697)))) severity failure;
    assert RAM(5698) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5698)))) severity failure;
    assert RAM(5699) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5699)))) severity failure;
    assert RAM(5700) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5700)))) severity failure;
    assert RAM(5701) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5701)))) severity failure;
    assert RAM(5702) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5702)))) severity failure;
    assert RAM(5703) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5703)))) severity failure;
    assert RAM(5704) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5704)))) severity failure;
    assert RAM(5705) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5705)))) severity failure;
    assert RAM(5706) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5706)))) severity failure;
    assert RAM(5707) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5707)))) severity failure;
    assert RAM(5708) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5708)))) severity failure;
    assert RAM(5709) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5709)))) severity failure;
    assert RAM(5710) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5710)))) severity failure;
    assert RAM(5711) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5711)))) severity failure;
    assert RAM(5712) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5712)))) severity failure;
    assert RAM(5713) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5713)))) severity failure;
    assert RAM(5714) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5714)))) severity failure;
    assert RAM(5715) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5715)))) severity failure;
    assert RAM(5716) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5716)))) severity failure;
    assert RAM(5717) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5717)))) severity failure;
    assert RAM(5718) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5718)))) severity failure;
    assert RAM(5719) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5719)))) severity failure;
    assert RAM(5720) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5720)))) severity failure;
    assert RAM(5721) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5721)))) severity failure;
    assert RAM(5722) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5722)))) severity failure;
    assert RAM(5723) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5723)))) severity failure;
    assert RAM(5724) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5724)))) severity failure;
    assert RAM(5725) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5725)))) severity failure;
    assert RAM(5726) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5726)))) severity failure;
    assert RAM(5727) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5727)))) severity failure;
    assert RAM(5728) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5728)))) severity failure;
    assert RAM(5729) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5729)))) severity failure;
    assert RAM(5730) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5730)))) severity failure;
    assert RAM(5731) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5731)))) severity failure;
    assert RAM(5732) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5732)))) severity failure;
    assert RAM(5733) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5733)))) severity failure;
    assert RAM(5734) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5734)))) severity failure;
    assert RAM(5735) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5735)))) severity failure;
    assert RAM(5736) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5736)))) severity failure;
    assert RAM(5737) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5737)))) severity failure;
    assert RAM(5738) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5738)))) severity failure;
    assert RAM(5739) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5739)))) severity failure;
    assert RAM(5740) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5740)))) severity failure;
    assert RAM(5741) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5741)))) severity failure;
    assert RAM(5742) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5742)))) severity failure;
    assert RAM(5743) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5743)))) severity failure;
    assert RAM(5744) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5744)))) severity failure;
    assert RAM(5745) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5745)))) severity failure;
    assert RAM(5746) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5746)))) severity failure;
    assert RAM(5747) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5747)))) severity failure;
    assert RAM(5748) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5748)))) severity failure;
    assert RAM(5749) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5749)))) severity failure;
    assert RAM(5750) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5750)))) severity failure;
    assert RAM(5751) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5751)))) severity failure;
    assert RAM(5752) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5752)))) severity failure;
    assert RAM(5753) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5753)))) severity failure;
    assert RAM(5754) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5754)))) severity failure;
    assert RAM(5755) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5755)))) severity failure;
    assert RAM(5756) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5756)))) severity failure;
    assert RAM(5757) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5757)))) severity failure;
    assert RAM(5758) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5758)))) severity failure;
    assert RAM(5759) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5759)))) severity failure;
    assert RAM(5760) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5760)))) severity failure;
    assert RAM(5761) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5761)))) severity failure;
    assert RAM(5762) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5762)))) severity failure;
    assert RAM(5763) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5763)))) severity failure;
    assert RAM(5764) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5764)))) severity failure;
    assert RAM(5765) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5765)))) severity failure;
    assert RAM(5766) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5766)))) severity failure;
    assert RAM(5767) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5767)))) severity failure;
    assert RAM(5768) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5768)))) severity failure;
    assert RAM(5769) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5769)))) severity failure;
    assert RAM(5770) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5770)))) severity failure;
    assert RAM(5771) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5771)))) severity failure;
    assert RAM(5772) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5772)))) severity failure;
    assert RAM(5773) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5773)))) severity failure;
    assert RAM(5774) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5774)))) severity failure;
    assert RAM(5775) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5775)))) severity failure;
    assert RAM(5776) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5776)))) severity failure;
    assert RAM(5777) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5777)))) severity failure;
    assert RAM(5778) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5778)))) severity failure;
    assert RAM(5779) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5779)))) severity failure;
    assert RAM(5780) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5780)))) severity failure;
    assert RAM(5781) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5781)))) severity failure;
    assert RAM(5782) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5782)))) severity failure;
    assert RAM(5783) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5783)))) severity failure;
    assert RAM(5784) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5784)))) severity failure;
    assert RAM(5785) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5785)))) severity failure;
    assert RAM(5786) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5786)))) severity failure;
    assert RAM(5787) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5787)))) severity failure;
    assert RAM(5788) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5788)))) severity failure;
    assert RAM(5789) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5789)))) severity failure;
    assert RAM(5790) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5790)))) severity failure;
    assert RAM(5791) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5791)))) severity failure;
    assert RAM(5792) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5792)))) severity failure;
    assert RAM(5793) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5793)))) severity failure;
    assert RAM(5794) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5794)))) severity failure;
    assert RAM(5795) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5795)))) severity failure;
    assert RAM(5796) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5796)))) severity failure;
    assert RAM(5797) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5797)))) severity failure;
    assert RAM(5798) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5798)))) severity failure;
    assert RAM(5799) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5799)))) severity failure;
    assert RAM(5800) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5800)))) severity failure;
    assert RAM(5801) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5801)))) severity failure;
    assert RAM(5802) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5802)))) severity failure;
    assert RAM(5803) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5803)))) severity failure;
    assert RAM(5804) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5804)))) severity failure;
    assert RAM(5805) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5805)))) severity failure;
    assert RAM(5806) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5806)))) severity failure;
    assert RAM(5807) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5807)))) severity failure;
    assert RAM(5808) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5808)))) severity failure;
    assert RAM(5809) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5809)))) severity failure;
    assert RAM(5810) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5810)))) severity failure;
    assert RAM(5811) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5811)))) severity failure;
    assert RAM(5812) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5812)))) severity failure;
    assert RAM(5813) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5813)))) severity failure;
    assert RAM(5814) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5814)))) severity failure;
    assert RAM(5815) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5815)))) severity failure;
    assert RAM(5816) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5816)))) severity failure;
    assert RAM(5817) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5817)))) severity failure;
    assert RAM(5818) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5818)))) severity failure;
    assert RAM(5819) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5819)))) severity failure;
    assert RAM(5820) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5820)))) severity failure;
    assert RAM(5821) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5821)))) severity failure;
    assert RAM(5822) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5822)))) severity failure;
    assert RAM(5823) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5823)))) severity failure;
    assert RAM(5824) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5824)))) severity failure;
    assert RAM(5825) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5825)))) severity failure;
    assert RAM(5826) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5826)))) severity failure;
    assert RAM(5827) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5827)))) severity failure;
    assert RAM(5828) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5828)))) severity failure;
    assert RAM(5829) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5829)))) severity failure;
    assert RAM(5830) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5830)))) severity failure;
    assert RAM(5831) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5831)))) severity failure;
    assert RAM(5832) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5832)))) severity failure;
    assert RAM(5833) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5833)))) severity failure;
    assert RAM(5834) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5834)))) severity failure;
    assert RAM(5835) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5835)))) severity failure;
    assert RAM(5836) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5836)))) severity failure;
    assert RAM(5837) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5837)))) severity failure;
    assert RAM(5838) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5838)))) severity failure;
    assert RAM(5839) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5839)))) severity failure;
    assert RAM(5840) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5840)))) severity failure;
    assert RAM(5841) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5841)))) severity failure;
    assert RAM(5842) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5842)))) severity failure;
    assert RAM(5843) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5843)))) severity failure;
    assert RAM(5844) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5844)))) severity failure;
    assert RAM(5845) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5845)))) severity failure;
    assert RAM(5846) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5846)))) severity failure;
    assert RAM(5847) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5847)))) severity failure;
    assert RAM(5848) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5848)))) severity failure;
    assert RAM(5849) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5849)))) severity failure;
    assert RAM(5850) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5850)))) severity failure;
    assert RAM(5851) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5851)))) severity failure;
    assert RAM(5852) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5852)))) severity failure;
    assert RAM(5853) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5853)))) severity failure;
    assert RAM(5854) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5854)))) severity failure;
    assert RAM(5855) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5855)))) severity failure;
    assert RAM(5856) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5856)))) severity failure;
    assert RAM(5857) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5857)))) severity failure;
    assert RAM(5858) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5858)))) severity failure;
    assert RAM(5859) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5859)))) severity failure;
    assert RAM(5860) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5860)))) severity failure;
    assert RAM(5861) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5861)))) severity failure;
    assert RAM(5862) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5862)))) severity failure;
    assert RAM(5863) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5863)))) severity failure;
    assert RAM(5864) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5864)))) severity failure;
    assert RAM(5865) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5865)))) severity failure;
    assert RAM(5866) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5866)))) severity failure;
    assert RAM(5867) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5867)))) severity failure;
    assert RAM(5868) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5868)))) severity failure;
    assert RAM(5869) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5869)))) severity failure;
    assert RAM(5870) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5870)))) severity failure;
    assert RAM(5871) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5871)))) severity failure;
    assert RAM(5872) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5872)))) severity failure;
    assert RAM(5873) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5873)))) severity failure;
    assert RAM(5874) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5874)))) severity failure;
    assert RAM(5875) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5875)))) severity failure;
    assert RAM(5876) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5876)))) severity failure;
    assert RAM(5877) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5877)))) severity failure;
    assert RAM(5878) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5878)))) severity failure;
    assert RAM(5879) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5879)))) severity failure;
    assert RAM(5880) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5880)))) severity failure;
    assert RAM(5881) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5881)))) severity failure;
    assert RAM(5882) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5882)))) severity failure;
    assert RAM(5883) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5883)))) severity failure;
    assert RAM(5884) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5884)))) severity failure;
    assert RAM(5885) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5885)))) severity failure;
    assert RAM(5886) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5886)))) severity failure;
    assert RAM(5887) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5887)))) severity failure;
    assert RAM(5888) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5888)))) severity failure;
    assert RAM(5889) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5889)))) severity failure;
    assert RAM(5890) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5890)))) severity failure;
    assert RAM(5891) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5891)))) severity failure;
    assert RAM(5892) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5892)))) severity failure;
    assert RAM(5893) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5893)))) severity failure;
    assert RAM(5894) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5894)))) severity failure;
    assert RAM(5895) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5895)))) severity failure;
    assert RAM(5896) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5896)))) severity failure;
    assert RAM(5897) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5897)))) severity failure;
    assert RAM(5898) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5898)))) severity failure;
    assert RAM(5899) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5899)))) severity failure;
    assert RAM(5900) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5900)))) severity failure;
    assert RAM(5901) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5901)))) severity failure;
    assert RAM(5902) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5902)))) severity failure;
    assert RAM(5903) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5903)))) severity failure;
    assert RAM(5904) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5904)))) severity failure;
    assert RAM(5905) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5905)))) severity failure;
    assert RAM(5906) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5906)))) severity failure;
    assert RAM(5907) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5907)))) severity failure;
    assert RAM(5908) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5908)))) severity failure;
    assert RAM(5909) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5909)))) severity failure;
    assert RAM(5910) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5910)))) severity failure;
    assert RAM(5911) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5911)))) severity failure;
    assert RAM(5912) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5912)))) severity failure;
    assert RAM(5913) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5913)))) severity failure;
    assert RAM(5914) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5914)))) severity failure;
    assert RAM(5915) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5915)))) severity failure;
    assert RAM(5916) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5916)))) severity failure;
    assert RAM(5917) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5917)))) severity failure;
    assert RAM(5918) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5918)))) severity failure;
    assert RAM(5919) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5919)))) severity failure;
    assert RAM(5920) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5920)))) severity failure;
    assert RAM(5921) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5921)))) severity failure;
    assert RAM(5922) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5922)))) severity failure;
    assert RAM(5923) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(5923)))) severity failure;
    assert RAM(5924) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5924)))) severity failure;
    assert RAM(5925) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5925)))) severity failure;
    assert RAM(5926) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5926)))) severity failure;
    assert RAM(5927) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5927)))) severity failure;
    assert RAM(5928) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5928)))) severity failure;
    assert RAM(5929) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5929)))) severity failure;
    assert RAM(5930) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5930)))) severity failure;
    assert RAM(5931) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5931)))) severity failure;
    assert RAM(5932) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(5932)))) severity failure;
    assert RAM(5933) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5933)))) severity failure;
    assert RAM(5934) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5934)))) severity failure;
    assert RAM(5935) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5935)))) severity failure;
    assert RAM(5936) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5936)))) severity failure;
    assert RAM(5937) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5937)))) severity failure;
    assert RAM(5938) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5938)))) severity failure;
    assert RAM(5939) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5939)))) severity failure;
    assert RAM(5940) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5940)))) severity failure;
    assert RAM(5941) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5941)))) severity failure;
    assert RAM(5942) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5942)))) severity failure;
    assert RAM(5943) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5943)))) severity failure;
    assert RAM(5944) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5944)))) severity failure;
    assert RAM(5945) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5945)))) severity failure;
    assert RAM(5946) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5946)))) severity failure;
    assert RAM(5947) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5947)))) severity failure;
    assert RAM(5948) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5948)))) severity failure;
    assert RAM(5949) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5949)))) severity failure;
    assert RAM(5950) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5950)))) severity failure;
    assert RAM(5951) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5951)))) severity failure;
    assert RAM(5952) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5952)))) severity failure;
    assert RAM(5953) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5953)))) severity failure;
    assert RAM(5954) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5954)))) severity failure;
    assert RAM(5955) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5955)))) severity failure;
    assert RAM(5956) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5956)))) severity failure;
    assert RAM(5957) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5957)))) severity failure;
    assert RAM(5958) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5958)))) severity failure;
    assert RAM(5959) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5959)))) severity failure;
    assert RAM(5960) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5960)))) severity failure;
    assert RAM(5961) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5961)))) severity failure;
    assert RAM(5962) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5962)))) severity failure;
    assert RAM(5963) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5963)))) severity failure;
    assert RAM(5964) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5964)))) severity failure;
    assert RAM(5965) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5965)))) severity failure;
    assert RAM(5966) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5966)))) severity failure;
    assert RAM(5967) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5967)))) severity failure;
    assert RAM(5968) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5968)))) severity failure;
    assert RAM(5969) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5969)))) severity failure;
    assert RAM(5970) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5970)))) severity failure;
    assert RAM(5971) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5971)))) severity failure;
    assert RAM(5972) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5972)))) severity failure;
    assert RAM(5973) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5973)))) severity failure;
    assert RAM(5974) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5974)))) severity failure;
    assert RAM(5975) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5975)))) severity failure;
    assert RAM(5976) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5976)))) severity failure;
    assert RAM(5977) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5977)))) severity failure;
    assert RAM(5978) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(5978)))) severity failure;
    assert RAM(5979) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5979)))) severity failure;
    assert RAM(5980) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(5980)))) severity failure;
    assert RAM(5981) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5981)))) severity failure;
    assert RAM(5982) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5982)))) severity failure;
    assert RAM(5983) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5983)))) severity failure;
    assert RAM(5984) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5984)))) severity failure;
    assert RAM(5985) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5985)))) severity failure;
    assert RAM(5986) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5986)))) severity failure;
    assert RAM(5987) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(5987)))) severity failure;
    assert RAM(5988) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5988)))) severity failure;
    assert RAM(5989) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5989)))) severity failure;
    assert RAM(5990) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5990)))) severity failure;
    assert RAM(5991) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5991)))) severity failure;
    assert RAM(5992) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5992)))) severity failure;
    assert RAM(5993) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(5993)))) severity failure;
    assert RAM(5994) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5994)))) severity failure;
    assert RAM(5995) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(5995)))) severity failure;
    assert RAM(5996) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5996)))) severity failure;
    assert RAM(5997) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5997)))) severity failure;
    assert RAM(5998) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(5998)))) severity failure;
    assert RAM(5999) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(5999)))) severity failure;
    assert RAM(6000) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6000)))) severity failure;
    assert RAM(6001) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6001)))) severity failure;
    assert RAM(6002) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6002)))) severity failure;
    assert RAM(6003) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6003)))) severity failure;
    assert RAM(6004) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6004)))) severity failure;
    assert RAM(6005) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6005)))) severity failure;
    assert RAM(6006) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6006)))) severity failure;
    assert RAM(6007) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6007)))) severity failure;
    assert RAM(6008) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6008)))) severity failure;
    assert RAM(6009) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6009)))) severity failure;
    assert RAM(6010) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6010)))) severity failure;
    assert RAM(6011) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6011)))) severity failure;
    assert RAM(6012) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6012)))) severity failure;
    assert RAM(6013) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6013)))) severity failure;
    assert RAM(6014) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6014)))) severity failure;
    assert RAM(6015) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6015)))) severity failure;
    assert RAM(6016) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6016)))) severity failure;
    assert RAM(6017) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6017)))) severity failure;
    assert RAM(6018) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6018)))) severity failure;
    assert RAM(6019) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6019)))) severity failure;
    assert RAM(6020) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6020)))) severity failure;
    assert RAM(6021) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6021)))) severity failure;
    assert RAM(6022) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6022)))) severity failure;
    assert RAM(6023) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6023)))) severity failure;
    assert RAM(6024) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6024)))) severity failure;
    assert RAM(6025) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6025)))) severity failure;
    assert RAM(6026) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6026)))) severity failure;
    assert RAM(6027) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6027)))) severity failure;
    assert RAM(6028) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6028)))) severity failure;
    assert RAM(6029) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6029)))) severity failure;
    assert RAM(6030) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6030)))) severity failure;
    assert RAM(6031) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6031)))) severity failure;
    assert RAM(6032) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6032)))) severity failure;
    assert RAM(6033) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6033)))) severity failure;
    assert RAM(6034) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6034)))) severity failure;
    assert RAM(6035) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6035)))) severity failure;
    assert RAM(6036) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6036)))) severity failure;
    assert RAM(6037) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6037)))) severity failure;
    assert RAM(6038) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6038)))) severity failure;
    assert RAM(6039) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6039)))) severity failure;
    assert RAM(6040) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6040)))) severity failure;
    assert RAM(6041) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6041)))) severity failure;
    assert RAM(6042) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6042)))) severity failure;
    assert RAM(6043) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6043)))) severity failure;
    assert RAM(6044) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6044)))) severity failure;
    assert RAM(6045) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6045)))) severity failure;
    assert RAM(6046) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6046)))) severity failure;
    assert RAM(6047) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6047)))) severity failure;
    assert RAM(6048) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6048)))) severity failure;
    assert RAM(6049) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6049)))) severity failure;
    assert RAM(6050) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6050)))) severity failure;
    assert RAM(6051) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6051)))) severity failure;
    assert RAM(6052) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6052)))) severity failure;
    assert RAM(6053) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6053)))) severity failure;
    assert RAM(6054) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6054)))) severity failure;
    assert RAM(6055) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6055)))) severity failure;
    assert RAM(6056) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6056)))) severity failure;
    assert RAM(6057) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6057)))) severity failure;
    assert RAM(6058) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6058)))) severity failure;
    assert RAM(6059) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6059)))) severity failure;
    assert RAM(6060) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6060)))) severity failure;
    assert RAM(6061) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6061)))) severity failure;
    assert RAM(6062) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6062)))) severity failure;
    assert RAM(6063) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6063)))) severity failure;
    assert RAM(6064) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6064)))) severity failure;
    assert RAM(6065) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6065)))) severity failure;
    assert RAM(6066) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6066)))) severity failure;
    assert RAM(6067) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6067)))) severity failure;
    assert RAM(6068) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6068)))) severity failure;
    assert RAM(6069) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6069)))) severity failure;
    assert RAM(6070) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6070)))) severity failure;
    assert RAM(6071) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6071)))) severity failure;
    assert RAM(6072) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6072)))) severity failure;
    assert RAM(6073) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6073)))) severity failure;
    assert RAM(6074) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6074)))) severity failure;
    assert RAM(6075) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6075)))) severity failure;
    assert RAM(6076) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6076)))) severity failure;
    assert RAM(6077) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6077)))) severity failure;
    assert RAM(6078) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6078)))) severity failure;
    assert RAM(6079) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6079)))) severity failure;
    assert RAM(6080) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6080)))) severity failure;
    assert RAM(6081) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6081)))) severity failure;
    assert RAM(6082) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6082)))) severity failure;
    assert RAM(6083) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6083)))) severity failure;
    assert RAM(6084) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6084)))) severity failure;
    assert RAM(6085) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6085)))) severity failure;
    assert RAM(6086) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6086)))) severity failure;
    assert RAM(6087) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6087)))) severity failure;
    assert RAM(6088) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6088)))) severity failure;
    assert RAM(6089) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6089)))) severity failure;
    assert RAM(6090) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6090)))) severity failure;
    assert RAM(6091) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6091)))) severity failure;
    assert RAM(6092) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6092)))) severity failure;
    assert RAM(6093) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6093)))) severity failure;
    assert RAM(6094) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6094)))) severity failure;
    assert RAM(6095) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6095)))) severity failure;
    assert RAM(6096) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6096)))) severity failure;
    assert RAM(6097) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6097)))) severity failure;
    assert RAM(6098) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6098)))) severity failure;
    assert RAM(6099) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6099)))) severity failure;
    assert RAM(6100) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6100)))) severity failure;
    assert RAM(6101) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6101)))) severity failure;
    assert RAM(6102) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6102)))) severity failure;
    assert RAM(6103) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6103)))) severity failure;
    assert RAM(6104) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6104)))) severity failure;
    assert RAM(6105) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6105)))) severity failure;
    assert RAM(6106) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6106)))) severity failure;
    assert RAM(6107) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6107)))) severity failure;
    assert RAM(6108) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6108)))) severity failure;
    assert RAM(6109) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6109)))) severity failure;
    assert RAM(6110) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6110)))) severity failure;
    assert RAM(6111) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6111)))) severity failure;
    assert RAM(6112) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6112)))) severity failure;
    assert RAM(6113) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6113)))) severity failure;
    assert RAM(6114) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6114)))) severity failure;
    assert RAM(6115) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6115)))) severity failure;
    assert RAM(6116) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6116)))) severity failure;
    assert RAM(6117) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6117)))) severity failure;
    assert RAM(6118) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6118)))) severity failure;
    assert RAM(6119) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6119)))) severity failure;
    assert RAM(6120) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6120)))) severity failure;
    assert RAM(6121) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6121)))) severity failure;
    assert RAM(6122) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6122)))) severity failure;
    assert RAM(6123) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6123)))) severity failure;
    assert RAM(6124) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6124)))) severity failure;
    assert RAM(6125) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6125)))) severity failure;
    assert RAM(6126) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6126)))) severity failure;
    assert RAM(6127) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6127)))) severity failure;
    assert RAM(6128) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6128)))) severity failure;
    assert RAM(6129) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6129)))) severity failure;
    assert RAM(6130) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6130)))) severity failure;
    assert RAM(6131) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6131)))) severity failure;
    assert RAM(6132) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6132)))) severity failure;
    assert RAM(6133) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6133)))) severity failure;
    assert RAM(6134) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6134)))) severity failure;
    assert RAM(6135) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6135)))) severity failure;
    assert RAM(6136) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6136)))) severity failure;
    assert RAM(6137) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6137)))) severity failure;
    assert RAM(6138) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6138)))) severity failure;
    assert RAM(6139) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6139)))) severity failure;
    assert RAM(6140) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6140)))) severity failure;
    assert RAM(6141) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6141)))) severity failure;
    assert RAM(6142) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6142)))) severity failure;
    assert RAM(6143) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6143)))) severity failure;
    assert RAM(6144) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6144)))) severity failure;
    assert RAM(6145) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6145)))) severity failure;
    assert RAM(6146) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6146)))) severity failure;
    assert RAM(6147) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6147)))) severity failure;
    assert RAM(6148) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6148)))) severity failure;
    assert RAM(6149) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6149)))) severity failure;
    assert RAM(6150) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6150)))) severity failure;
    assert RAM(6151) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6151)))) severity failure;
    assert RAM(6152) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6152)))) severity failure;
    assert RAM(6153) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6153)))) severity failure;
    assert RAM(6154) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6154)))) severity failure;
    assert RAM(6155) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6155)))) severity failure;
    assert RAM(6156) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6156)))) severity failure;
    assert RAM(6157) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6157)))) severity failure;
    assert RAM(6158) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6158)))) severity failure;
    assert RAM(6159) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6159)))) severity failure;
    assert RAM(6160) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6160)))) severity failure;
    assert RAM(6161) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6161)))) severity failure;
    assert RAM(6162) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6162)))) severity failure;
    assert RAM(6163) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6163)))) severity failure;
    assert RAM(6164) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6164)))) severity failure;
    assert RAM(6165) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6165)))) severity failure;
    assert RAM(6166) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6166)))) severity failure;
    assert RAM(6167) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6167)))) severity failure;
    assert RAM(6168) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6168)))) severity failure;
    assert RAM(6169) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6169)))) severity failure;
    assert RAM(6170) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6170)))) severity failure;
    assert RAM(6171) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6171)))) severity failure;
    assert RAM(6172) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6172)))) severity failure;
    assert RAM(6173) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6173)))) severity failure;
    assert RAM(6174) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6174)))) severity failure;
    assert RAM(6175) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6175)))) severity failure;
    assert RAM(6176) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6176)))) severity failure;
    assert RAM(6177) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6177)))) severity failure;
    assert RAM(6178) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6178)))) severity failure;
    assert RAM(6179) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6179)))) severity failure;
    assert RAM(6180) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6180)))) severity failure;
    assert RAM(6181) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6181)))) severity failure;
    assert RAM(6182) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6182)))) severity failure;
    assert RAM(6183) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6183)))) severity failure;
    assert RAM(6184) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6184)))) severity failure;
    assert RAM(6185) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6185)))) severity failure;
    assert RAM(6186) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6186)))) severity failure;
    assert RAM(6187) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6187)))) severity failure;
    assert RAM(6188) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6188)))) severity failure;
    assert RAM(6189) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6189)))) severity failure;
    assert RAM(6190) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6190)))) severity failure;
    assert RAM(6191) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6191)))) severity failure;
    assert RAM(6192) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6192)))) severity failure;
    assert RAM(6193) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6193)))) severity failure;
    assert RAM(6194) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6194)))) severity failure;
    assert RAM(6195) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6195)))) severity failure;
    assert RAM(6196) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6196)))) severity failure;
    assert RAM(6197) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6197)))) severity failure;
    assert RAM(6198) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6198)))) severity failure;
    assert RAM(6199) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6199)))) severity failure;
    assert RAM(6200) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6200)))) severity failure;
    assert RAM(6201) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6201)))) severity failure;
    assert RAM(6202) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6202)))) severity failure;
    assert RAM(6203) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6203)))) severity failure;
    assert RAM(6204) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6204)))) severity failure;
    assert RAM(6205) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6205)))) severity failure;
    assert RAM(6206) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6206)))) severity failure;
    assert RAM(6207) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6207)))) severity failure;
    assert RAM(6208) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6208)))) severity failure;
    assert RAM(6209) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6209)))) severity failure;
    assert RAM(6210) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6210)))) severity failure;
    assert RAM(6211) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6211)))) severity failure;
    assert RAM(6212) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6212)))) severity failure;
    assert RAM(6213) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6213)))) severity failure;
    assert RAM(6214) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6214)))) severity failure;
    assert RAM(6215) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6215)))) severity failure;
    assert RAM(6216) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6216)))) severity failure;
    assert RAM(6217) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6217)))) severity failure;
    assert RAM(6218) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6218)))) severity failure;
    assert RAM(6219) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6219)))) severity failure;
    assert RAM(6220) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6220)))) severity failure;
    assert RAM(6221) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6221)))) severity failure;
    assert RAM(6222) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6222)))) severity failure;
    assert RAM(6223) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6223)))) severity failure;
    assert RAM(6224) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6224)))) severity failure;
    assert RAM(6225) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6225)))) severity failure;
    assert RAM(6226) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6226)))) severity failure;
    assert RAM(6227) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6227)))) severity failure;
    assert RAM(6228) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6228)))) severity failure;
    assert RAM(6229) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6229)))) severity failure;
    assert RAM(6230) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6230)))) severity failure;
    assert RAM(6231) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6231)))) severity failure;
    assert RAM(6232) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6232)))) severity failure;
    assert RAM(6233) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6233)))) severity failure;
    assert RAM(6234) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6234)))) severity failure;
    assert RAM(6235) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6235)))) severity failure;
    assert RAM(6236) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6236)))) severity failure;
    assert RAM(6237) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6237)))) severity failure;
    assert RAM(6238) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6238)))) severity failure;
    assert RAM(6239) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6239)))) severity failure;
    assert RAM(6240) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6240)))) severity failure;
    assert RAM(6241) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6241)))) severity failure;
    assert RAM(6242) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6242)))) severity failure;
    assert RAM(6243) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6243)))) severity failure;
    assert RAM(6244) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6244)))) severity failure;
    assert RAM(6245) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6245)))) severity failure;
    assert RAM(6246) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6246)))) severity failure;
    assert RAM(6247) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6247)))) severity failure;
    assert RAM(6248) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6248)))) severity failure;
    assert RAM(6249) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6249)))) severity failure;
    assert RAM(6250) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6250)))) severity failure;
    assert RAM(6251) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6251)))) severity failure;
    assert RAM(6252) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6252)))) severity failure;
    assert RAM(6253) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6253)))) severity failure;
    assert RAM(6254) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6254)))) severity failure;
    assert RAM(6255) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6255)))) severity failure;
    assert RAM(6256) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6256)))) severity failure;
    assert RAM(6257) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6257)))) severity failure;
    assert RAM(6258) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6258)))) severity failure;
    assert RAM(6259) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6259)))) severity failure;
    assert RAM(6260) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6260)))) severity failure;
    assert RAM(6261) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6261)))) severity failure;
    assert RAM(6262) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6262)))) severity failure;
    assert RAM(6263) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6263)))) severity failure;
    assert RAM(6264) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6264)))) severity failure;
    assert RAM(6265) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6265)))) severity failure;
    assert RAM(6266) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6266)))) severity failure;
    assert RAM(6267) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6267)))) severity failure;
    assert RAM(6268) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6268)))) severity failure;
    assert RAM(6269) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6269)))) severity failure;
    assert RAM(6270) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6270)))) severity failure;
    assert RAM(6271) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6271)))) severity failure;
    assert RAM(6272) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6272)))) severity failure;
    assert RAM(6273) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6273)))) severity failure;
    assert RAM(6274) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6274)))) severity failure;
    assert RAM(6275) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6275)))) severity failure;
    assert RAM(6276) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6276)))) severity failure;
    assert RAM(6277) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6277)))) severity failure;
    assert RAM(6278) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6278)))) severity failure;
    assert RAM(6279) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6279)))) severity failure;
    assert RAM(6280) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6280)))) severity failure;
    assert RAM(6281) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6281)))) severity failure;
    assert RAM(6282) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6282)))) severity failure;
    assert RAM(6283) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6283)))) severity failure;
    assert RAM(6284) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6284)))) severity failure;
    assert RAM(6285) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6285)))) severity failure;
    assert RAM(6286) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6286)))) severity failure;
    assert RAM(6287) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6287)))) severity failure;
    assert RAM(6288) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6288)))) severity failure;
    assert RAM(6289) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6289)))) severity failure;
    assert RAM(6290) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6290)))) severity failure;
    assert RAM(6291) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6291)))) severity failure;
    assert RAM(6292) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6292)))) severity failure;
    assert RAM(6293) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6293)))) severity failure;
    assert RAM(6294) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6294)))) severity failure;
    assert RAM(6295) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6295)))) severity failure;
    assert RAM(6296) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6296)))) severity failure;
    assert RAM(6297) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6297)))) severity failure;
    assert RAM(6298) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6298)))) severity failure;
    assert RAM(6299) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6299)))) severity failure;
    assert RAM(6300) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6300)))) severity failure;
    assert RAM(6301) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6301)))) severity failure;
    assert RAM(6302) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6302)))) severity failure;
    assert RAM(6303) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6303)))) severity failure;
    assert RAM(6304) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6304)))) severity failure;
    assert RAM(6305) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6305)))) severity failure;
    assert RAM(6306) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6306)))) severity failure;
    assert RAM(6307) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6307)))) severity failure;
    assert RAM(6308) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6308)))) severity failure;
    assert RAM(6309) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6309)))) severity failure;
    assert RAM(6310) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6310)))) severity failure;
    assert RAM(6311) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6311)))) severity failure;
    assert RAM(6312) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6312)))) severity failure;
    assert RAM(6313) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6313)))) severity failure;
    assert RAM(6314) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6314)))) severity failure;
    assert RAM(6315) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6315)))) severity failure;
    assert RAM(6316) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6316)))) severity failure;
    assert RAM(6317) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6317)))) severity failure;
    assert RAM(6318) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6318)))) severity failure;
    assert RAM(6319) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6319)))) severity failure;
    assert RAM(6320) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6320)))) severity failure;
    assert RAM(6321) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6321)))) severity failure;
    assert RAM(6322) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6322)))) severity failure;
    assert RAM(6323) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6323)))) severity failure;
    assert RAM(6324) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6324)))) severity failure;
    assert RAM(6325) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6325)))) severity failure;
    assert RAM(6326) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6326)))) severity failure;
    assert RAM(6327) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6327)))) severity failure;
    assert RAM(6328) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6328)))) severity failure;
    assert RAM(6329) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6329)))) severity failure;
    assert RAM(6330) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6330)))) severity failure;
    assert RAM(6331) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6331)))) severity failure;
    assert RAM(6332) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6332)))) severity failure;
    assert RAM(6333) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6333)))) severity failure;
    assert RAM(6334) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6334)))) severity failure;
    assert RAM(6335) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6335)))) severity failure;
    assert RAM(6336) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6336)))) severity failure;
    assert RAM(6337) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6337)))) severity failure;
    assert RAM(6338) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6338)))) severity failure;
    assert RAM(6339) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6339)))) severity failure;
    assert RAM(6340) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6340)))) severity failure;
    assert RAM(6341) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6341)))) severity failure;
    assert RAM(6342) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6342)))) severity failure;
    assert RAM(6343) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6343)))) severity failure;
    assert RAM(6344) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6344)))) severity failure;
    assert RAM(6345) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6345)))) severity failure;
    assert RAM(6346) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6346)))) severity failure;
    assert RAM(6347) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6347)))) severity failure;
    assert RAM(6348) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6348)))) severity failure;
    assert RAM(6349) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6349)))) severity failure;
    assert RAM(6350) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6350)))) severity failure;
    assert RAM(6351) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6351)))) severity failure;
    assert RAM(6352) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6352)))) severity failure;
    assert RAM(6353) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6353)))) severity failure;
    assert RAM(6354) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6354)))) severity failure;
    assert RAM(6355) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6355)))) severity failure;
    assert RAM(6356) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6356)))) severity failure;
    assert RAM(6357) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6357)))) severity failure;
    assert RAM(6358) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6358)))) severity failure;
    assert RAM(6359) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6359)))) severity failure;
    assert RAM(6360) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6360)))) severity failure;
    assert RAM(6361) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6361)))) severity failure;
    assert RAM(6362) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6362)))) severity failure;
    assert RAM(6363) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6363)))) severity failure;
    assert RAM(6364) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6364)))) severity failure;
    assert RAM(6365) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6365)))) severity failure;
    assert RAM(6366) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6366)))) severity failure;
    assert RAM(6367) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6367)))) severity failure;
    assert RAM(6368) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6368)))) severity failure;
    assert RAM(6369) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6369)))) severity failure;
    assert RAM(6370) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6370)))) severity failure;
    assert RAM(6371) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6371)))) severity failure;
    assert RAM(6372) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6372)))) severity failure;
    assert RAM(6373) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6373)))) severity failure;
    assert RAM(6374) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6374)))) severity failure;
    assert RAM(6375) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6375)))) severity failure;
    assert RAM(6376) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6376)))) severity failure;
    assert RAM(6377) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6377)))) severity failure;
    assert RAM(6378) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6378)))) severity failure;
    assert RAM(6379) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6379)))) severity failure;
    assert RAM(6380) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6380)))) severity failure;
    assert RAM(6381) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6381)))) severity failure;
    assert RAM(6382) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6382)))) severity failure;
    assert RAM(6383) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6383)))) severity failure;
    assert RAM(6384) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6384)))) severity failure;
    assert RAM(6385) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6385)))) severity failure;
    assert RAM(6386) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6386)))) severity failure;
    assert RAM(6387) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6387)))) severity failure;
    assert RAM(6388) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6388)))) severity failure;
    assert RAM(6389) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6389)))) severity failure;
    assert RAM(6390) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6390)))) severity failure;
    assert RAM(6391) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6391)))) severity failure;
    assert RAM(6392) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6392)))) severity failure;
    assert RAM(6393) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6393)))) severity failure;
    assert RAM(6394) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6394)))) severity failure;
    assert RAM(6395) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6395)))) severity failure;
    assert RAM(6396) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6396)))) severity failure;
    assert RAM(6397) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6397)))) severity failure;
    assert RAM(6398) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6398)))) severity failure;
    assert RAM(6399) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6399)))) severity failure;
    assert RAM(6400) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6400)))) severity failure;
    assert RAM(6401) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6401)))) severity failure;
    assert RAM(6402) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6402)))) severity failure;
    assert RAM(6403) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6403)))) severity failure;
    assert RAM(6404) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6404)))) severity failure;
    assert RAM(6405) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6405)))) severity failure;
    assert RAM(6406) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6406)))) severity failure;
    assert RAM(6407) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6407)))) severity failure;
    assert RAM(6408) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6408)))) severity failure;
    assert RAM(6409) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6409)))) severity failure;
    assert RAM(6410) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6410)))) severity failure;
    assert RAM(6411) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6411)))) severity failure;
    assert RAM(6412) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6412)))) severity failure;
    assert RAM(6413) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6413)))) severity failure;
    assert RAM(6414) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6414)))) severity failure;
    assert RAM(6415) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6415)))) severity failure;
    assert RAM(6416) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6416)))) severity failure;
    assert RAM(6417) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6417)))) severity failure;
    assert RAM(6418) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6418)))) severity failure;
    assert RAM(6419) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6419)))) severity failure;
    assert RAM(6420) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6420)))) severity failure;
    assert RAM(6421) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6421)))) severity failure;
    assert RAM(6422) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6422)))) severity failure;
    assert RAM(6423) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6423)))) severity failure;
    assert RAM(6424) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6424)))) severity failure;
    assert RAM(6425) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6425)))) severity failure;
    assert RAM(6426) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6426)))) severity failure;
    assert RAM(6427) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6427)))) severity failure;
    assert RAM(6428) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6428)))) severity failure;
    assert RAM(6429) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6429)))) severity failure;
    assert RAM(6430) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6430)))) severity failure;
    assert RAM(6431) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6431)))) severity failure;
    assert RAM(6432) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6432)))) severity failure;
    assert RAM(6433) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6433)))) severity failure;
    assert RAM(6434) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6434)))) severity failure;
    assert RAM(6435) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6435)))) severity failure;
    assert RAM(6436) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6436)))) severity failure;
    assert RAM(6437) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6437)))) severity failure;
    assert RAM(6438) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6438)))) severity failure;
    assert RAM(6439) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6439)))) severity failure;
    assert RAM(6440) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6440)))) severity failure;
    assert RAM(6441) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6441)))) severity failure;
    assert RAM(6442) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6442)))) severity failure;
    assert RAM(6443) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6443)))) severity failure;
    assert RAM(6444) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6444)))) severity failure;
    assert RAM(6445) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6445)))) severity failure;
    assert RAM(6446) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6446)))) severity failure;
    assert RAM(6447) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6447)))) severity failure;
    assert RAM(6448) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6448)))) severity failure;
    assert RAM(6449) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6449)))) severity failure;
    assert RAM(6450) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6450)))) severity failure;
    assert RAM(6451) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6451)))) severity failure;
    assert RAM(6452) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6452)))) severity failure;
    assert RAM(6453) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6453)))) severity failure;
    assert RAM(6454) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6454)))) severity failure;
    assert RAM(6455) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6455)))) severity failure;
    assert RAM(6456) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6456)))) severity failure;
    assert RAM(6457) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6457)))) severity failure;
    assert RAM(6458) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6458)))) severity failure;
    assert RAM(6459) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6459)))) severity failure;
    assert RAM(6460) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6460)))) severity failure;
    assert RAM(6461) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6461)))) severity failure;
    assert RAM(6462) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6462)))) severity failure;
    assert RAM(6463) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6463)))) severity failure;
    assert RAM(6464) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6464)))) severity failure;
    assert RAM(6465) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6465)))) severity failure;
    assert RAM(6466) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6466)))) severity failure;
    assert RAM(6467) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6467)))) severity failure;
    assert RAM(6468) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6468)))) severity failure;
    assert RAM(6469) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6469)))) severity failure;
    assert RAM(6470) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6470)))) severity failure;
    assert RAM(6471) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6471)))) severity failure;
    assert RAM(6472) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6472)))) severity failure;
    assert RAM(6473) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6473)))) severity failure;
    assert RAM(6474) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6474)))) severity failure;
    assert RAM(6475) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6475)))) severity failure;
    assert RAM(6476) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6476)))) severity failure;
    assert RAM(6477) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6477)))) severity failure;
    assert RAM(6478) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6478)))) severity failure;
    assert RAM(6479) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6479)))) severity failure;
    assert RAM(6480) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6480)))) severity failure;
    assert RAM(6481) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6481)))) severity failure;
    assert RAM(6482) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6482)))) severity failure;
    assert RAM(6483) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6483)))) severity failure;
    assert RAM(6484) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6484)))) severity failure;
    assert RAM(6485) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6485)))) severity failure;
    assert RAM(6486) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6486)))) severity failure;
    assert RAM(6487) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6487)))) severity failure;
    assert RAM(6488) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6488)))) severity failure;
    assert RAM(6489) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6489)))) severity failure;
    assert RAM(6490) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6490)))) severity failure;
    assert RAM(6491) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6491)))) severity failure;
    assert RAM(6492) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6492)))) severity failure;
    assert RAM(6493) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6493)))) severity failure;
    assert RAM(6494) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6494)))) severity failure;
    assert RAM(6495) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6495)))) severity failure;
    assert RAM(6496) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6496)))) severity failure;
    assert RAM(6497) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6497)))) severity failure;
    assert RAM(6498) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6498)))) severity failure;
    assert RAM(6499) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6499)))) severity failure;
    assert RAM(6500) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6500)))) severity failure;
    assert RAM(6501) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6501)))) severity failure;
    assert RAM(6502) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6502)))) severity failure;
    assert RAM(6503) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6503)))) severity failure;
    assert RAM(6504) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6504)))) severity failure;
    assert RAM(6505) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6505)))) severity failure;
    assert RAM(6506) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6506)))) severity failure;
    assert RAM(6507) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6507)))) severity failure;
    assert RAM(6508) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6508)))) severity failure;
    assert RAM(6509) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6509)))) severity failure;
    assert RAM(6510) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6510)))) severity failure;
    assert RAM(6511) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6511)))) severity failure;
    assert RAM(6512) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6512)))) severity failure;
    assert RAM(6513) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6513)))) severity failure;
    assert RAM(6514) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6514)))) severity failure;
    assert RAM(6515) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6515)))) severity failure;
    assert RAM(6516) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6516)))) severity failure;
    assert RAM(6517) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6517)))) severity failure;
    assert RAM(6518) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6518)))) severity failure;
    assert RAM(6519) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6519)))) severity failure;
    assert RAM(6520) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6520)))) severity failure;
    assert RAM(6521) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6521)))) severity failure;
    assert RAM(6522) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6522)))) severity failure;
    assert RAM(6523) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6523)))) severity failure;
    assert RAM(6524) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6524)))) severity failure;
    assert RAM(6525) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6525)))) severity failure;
    assert RAM(6526) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6526)))) severity failure;
    assert RAM(6527) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6527)))) severity failure;
    assert RAM(6528) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6528)))) severity failure;
    assert RAM(6529) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6529)))) severity failure;
    assert RAM(6530) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6530)))) severity failure;
    assert RAM(6531) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6531)))) severity failure;
    assert RAM(6532) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6532)))) severity failure;
    assert RAM(6533) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6533)))) severity failure;
    assert RAM(6534) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6534)))) severity failure;
    assert RAM(6535) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6535)))) severity failure;
    assert RAM(6536) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6536)))) severity failure;
    assert RAM(6537) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6537)))) severity failure;
    assert RAM(6538) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6538)))) severity failure;
    assert RAM(6539) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6539)))) severity failure;
    assert RAM(6540) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6540)))) severity failure;
    assert RAM(6541) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6541)))) severity failure;
    assert RAM(6542) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6542)))) severity failure;
    assert RAM(6543) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6543)))) severity failure;
    assert RAM(6544) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6544)))) severity failure;
    assert RAM(6545) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6545)))) severity failure;
    assert RAM(6546) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6546)))) severity failure;
    assert RAM(6547) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6547)))) severity failure;
    assert RAM(6548) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6548)))) severity failure;
    assert RAM(6549) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6549)))) severity failure;
    assert RAM(6550) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6550)))) severity failure;
    assert RAM(6551) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6551)))) severity failure;
    assert RAM(6552) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6552)))) severity failure;
    assert RAM(6553) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6553)))) severity failure;
    assert RAM(6554) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6554)))) severity failure;
    assert RAM(6555) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6555)))) severity failure;
    assert RAM(6556) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6556)))) severity failure;
    assert RAM(6557) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6557)))) severity failure;
    assert RAM(6558) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6558)))) severity failure;
    assert RAM(6559) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6559)))) severity failure;
    assert RAM(6560) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6560)))) severity failure;
    assert RAM(6561) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6561)))) severity failure;
    assert RAM(6562) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6562)))) severity failure;
    assert RAM(6563) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6563)))) severity failure;
    assert RAM(6564) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6564)))) severity failure;
    assert RAM(6565) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6565)))) severity failure;
    assert RAM(6566) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6566)))) severity failure;
    assert RAM(6567) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6567)))) severity failure;
    assert RAM(6568) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6568)))) severity failure;
    assert RAM(6569) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6569)))) severity failure;
    assert RAM(6570) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6570)))) severity failure;
    assert RAM(6571) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6571)))) severity failure;
    assert RAM(6572) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6572)))) severity failure;
    assert RAM(6573) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6573)))) severity failure;
    assert RAM(6574) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6574)))) severity failure;
    assert RAM(6575) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6575)))) severity failure;
    assert RAM(6576) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6576)))) severity failure;
    assert RAM(6577) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6577)))) severity failure;
    assert RAM(6578) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6578)))) severity failure;
    assert RAM(6579) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6579)))) severity failure;
    assert RAM(6580) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6580)))) severity failure;
    assert RAM(6581) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6581)))) severity failure;
    assert RAM(6582) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6582)))) severity failure;
    assert RAM(6583) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6583)))) severity failure;
    assert RAM(6584) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6584)))) severity failure;
    assert RAM(6585) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6585)))) severity failure;
    assert RAM(6586) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6586)))) severity failure;
    assert RAM(6587) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6587)))) severity failure;
    assert RAM(6588) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6588)))) severity failure;
    assert RAM(6589) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6589)))) severity failure;
    assert RAM(6590) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6590)))) severity failure;
    assert RAM(6591) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6591)))) severity failure;
    assert RAM(6592) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6592)))) severity failure;
    assert RAM(6593) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6593)))) severity failure;
    assert RAM(6594) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6594)))) severity failure;
    assert RAM(6595) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6595)))) severity failure;
    assert RAM(6596) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6596)))) severity failure;
    assert RAM(6597) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6597)))) severity failure;
    assert RAM(6598) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6598)))) severity failure;
    assert RAM(6599) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6599)))) severity failure;
    assert RAM(6600) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6600)))) severity failure;
    assert RAM(6601) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6601)))) severity failure;
    assert RAM(6602) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6602)))) severity failure;
    assert RAM(6603) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6603)))) severity failure;
    assert RAM(6604) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6604)))) severity failure;
    assert RAM(6605) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6605)))) severity failure;
    assert RAM(6606) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6606)))) severity failure;
    assert RAM(6607) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6607)))) severity failure;
    assert RAM(6608) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6608)))) severity failure;
    assert RAM(6609) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6609)))) severity failure;
    assert RAM(6610) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6610)))) severity failure;
    assert RAM(6611) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6611)))) severity failure;
    assert RAM(6612) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6612)))) severity failure;
    assert RAM(6613) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6613)))) severity failure;
    assert RAM(6614) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6614)))) severity failure;
    assert RAM(6615) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6615)))) severity failure;
    assert RAM(6616) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6616)))) severity failure;
    assert RAM(6617) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6617)))) severity failure;
    assert RAM(6618) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6618)))) severity failure;
    assert RAM(6619) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6619)))) severity failure;
    assert RAM(6620) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6620)))) severity failure;
    assert RAM(6621) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6621)))) severity failure;
    assert RAM(6622) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6622)))) severity failure;
    assert RAM(6623) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6623)))) severity failure;
    assert RAM(6624) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6624)))) severity failure;
    assert RAM(6625) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6625)))) severity failure;
    assert RAM(6626) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6626)))) severity failure;
    assert RAM(6627) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6627)))) severity failure;
    assert RAM(6628) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6628)))) severity failure;
    assert RAM(6629) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6629)))) severity failure;
    assert RAM(6630) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6630)))) severity failure;
    assert RAM(6631) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6631)))) severity failure;
    assert RAM(6632) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6632)))) severity failure;
    assert RAM(6633) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6633)))) severity failure;
    assert RAM(6634) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6634)))) severity failure;
    assert RAM(6635) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6635)))) severity failure;
    assert RAM(6636) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6636)))) severity failure;
    assert RAM(6637) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6637)))) severity failure;
    assert RAM(6638) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6638)))) severity failure;
    assert RAM(6639) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6639)))) severity failure;
    assert RAM(6640) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6640)))) severity failure;
    assert RAM(6641) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6641)))) severity failure;
    assert RAM(6642) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6642)))) severity failure;
    assert RAM(6643) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6643)))) severity failure;
    assert RAM(6644) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6644)))) severity failure;
    assert RAM(6645) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6645)))) severity failure;
    assert RAM(6646) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6646)))) severity failure;
    assert RAM(6647) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6647)))) severity failure;
    assert RAM(6648) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6648)))) severity failure;
    assert RAM(6649) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6649)))) severity failure;
    assert RAM(6650) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6650)))) severity failure;
    assert RAM(6651) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6651)))) severity failure;
    assert RAM(6652) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6652)))) severity failure;
    assert RAM(6653) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6653)))) severity failure;
    assert RAM(6654) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6654)))) severity failure;
    assert RAM(6655) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6655)))) severity failure;
    assert RAM(6656) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6656)))) severity failure;
    assert RAM(6657) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6657)))) severity failure;
    assert RAM(6658) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6658)))) severity failure;
    assert RAM(6659) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6659)))) severity failure;
    assert RAM(6660) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6660)))) severity failure;
    assert RAM(6661) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6661)))) severity failure;
    assert RAM(6662) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6662)))) severity failure;
    assert RAM(6663) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6663)))) severity failure;
    assert RAM(6664) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6664)))) severity failure;
    assert RAM(6665) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6665)))) severity failure;
    assert RAM(6666) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6666)))) severity failure;
    assert RAM(6667) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6667)))) severity failure;
    assert RAM(6668) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6668)))) severity failure;
    assert RAM(6669) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6669)))) severity failure;
    assert RAM(6670) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6670)))) severity failure;
    assert RAM(6671) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6671)))) severity failure;
    assert RAM(6672) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6672)))) severity failure;
    assert RAM(6673) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6673)))) severity failure;
    assert RAM(6674) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6674)))) severity failure;
    assert RAM(6675) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6675)))) severity failure;
    assert RAM(6676) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6676)))) severity failure;
    assert RAM(6677) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6677)))) severity failure;
    assert RAM(6678) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6678)))) severity failure;
    assert RAM(6679) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6679)))) severity failure;
    assert RAM(6680) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6680)))) severity failure;
    assert RAM(6681) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6681)))) severity failure;
    assert RAM(6682) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6682)))) severity failure;
    assert RAM(6683) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6683)))) severity failure;
    assert RAM(6684) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6684)))) severity failure;
    assert RAM(6685) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6685)))) severity failure;
    assert RAM(6686) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6686)))) severity failure;
    assert RAM(6687) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6687)))) severity failure;
    assert RAM(6688) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6688)))) severity failure;
    assert RAM(6689) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6689)))) severity failure;
    assert RAM(6690) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6690)))) severity failure;
    assert RAM(6691) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6691)))) severity failure;
    assert RAM(6692) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6692)))) severity failure;
    assert RAM(6693) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6693)))) severity failure;
    assert RAM(6694) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6694)))) severity failure;
    assert RAM(6695) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6695)))) severity failure;
    assert RAM(6696) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6696)))) severity failure;
    assert RAM(6697) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6697)))) severity failure;
    assert RAM(6698) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6698)))) severity failure;
    assert RAM(6699) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6699)))) severity failure;
    assert RAM(6700) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6700)))) severity failure;
    assert RAM(6701) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6701)))) severity failure;
    assert RAM(6702) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6702)))) severity failure;
    assert RAM(6703) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6703)))) severity failure;
    assert RAM(6704) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6704)))) severity failure;
    assert RAM(6705) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6705)))) severity failure;
    assert RAM(6706) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6706)))) severity failure;
    assert RAM(6707) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6707)))) severity failure;
    assert RAM(6708) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6708)))) severity failure;
    assert RAM(6709) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6709)))) severity failure;
    assert RAM(6710) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6710)))) severity failure;
    assert RAM(6711) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6711)))) severity failure;
    assert RAM(6712) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6712)))) severity failure;
    assert RAM(6713) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6713)))) severity failure;
    assert RAM(6714) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6714)))) severity failure;
    assert RAM(6715) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6715)))) severity failure;
    assert RAM(6716) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6716)))) severity failure;
    assert RAM(6717) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6717)))) severity failure;
    assert RAM(6718) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6718)))) severity failure;
    assert RAM(6719) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6719)))) severity failure;
    assert RAM(6720) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6720)))) severity failure;
    assert RAM(6721) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6721)))) severity failure;
    assert RAM(6722) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6722)))) severity failure;
    assert RAM(6723) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6723)))) severity failure;
    assert RAM(6724) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6724)))) severity failure;
    assert RAM(6725) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6725)))) severity failure;
    assert RAM(6726) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6726)))) severity failure;
    assert RAM(6727) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6727)))) severity failure;
    assert RAM(6728) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6728)))) severity failure;
    assert RAM(6729) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6729)))) severity failure;
    assert RAM(6730) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6730)))) severity failure;
    assert RAM(6731) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6731)))) severity failure;
    assert RAM(6732) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6732)))) severity failure;
    assert RAM(6733) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6733)))) severity failure;
    assert RAM(6734) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6734)))) severity failure;
    assert RAM(6735) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6735)))) severity failure;
    assert RAM(6736) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6736)))) severity failure;
    assert RAM(6737) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6737)))) severity failure;
    assert RAM(6738) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6738)))) severity failure;
    assert RAM(6739) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6739)))) severity failure;
    assert RAM(6740) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6740)))) severity failure;
    assert RAM(6741) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6741)))) severity failure;
    assert RAM(6742) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6742)))) severity failure;
    assert RAM(6743) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6743)))) severity failure;
    assert RAM(6744) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6744)))) severity failure;
    assert RAM(6745) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6745)))) severity failure;
    assert RAM(6746) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6746)))) severity failure;
    assert RAM(6747) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6747)))) severity failure;
    assert RAM(6748) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6748)))) severity failure;
    assert RAM(6749) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6749)))) severity failure;
    assert RAM(6750) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6750)))) severity failure;
    assert RAM(6751) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6751)))) severity failure;
    assert RAM(6752) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6752)))) severity failure;
    assert RAM(6753) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6753)))) severity failure;
    assert RAM(6754) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6754)))) severity failure;
    assert RAM(6755) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6755)))) severity failure;
    assert RAM(6756) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6756)))) severity failure;
    assert RAM(6757) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6757)))) severity failure;
    assert RAM(6758) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6758)))) severity failure;
    assert RAM(6759) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6759)))) severity failure;
    assert RAM(6760) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6760)))) severity failure;
    assert RAM(6761) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6761)))) severity failure;
    assert RAM(6762) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6762)))) severity failure;
    assert RAM(6763) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6763)))) severity failure;
    assert RAM(6764) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6764)))) severity failure;
    assert RAM(6765) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6765)))) severity failure;
    assert RAM(6766) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6766)))) severity failure;
    assert RAM(6767) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6767)))) severity failure;
    assert RAM(6768) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6768)))) severity failure;
    assert RAM(6769) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6769)))) severity failure;
    assert RAM(6770) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6770)))) severity failure;
    assert RAM(6771) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6771)))) severity failure;
    assert RAM(6772) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6772)))) severity failure;
    assert RAM(6773) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6773)))) severity failure;
    assert RAM(6774) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6774)))) severity failure;
    assert RAM(6775) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6775)))) severity failure;
    assert RAM(6776) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6776)))) severity failure;
    assert RAM(6777) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6777)))) severity failure;
    assert RAM(6778) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6778)))) severity failure;
    assert RAM(6779) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6779)))) severity failure;
    assert RAM(6780) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6780)))) severity failure;
    assert RAM(6781) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6781)))) severity failure;
    assert RAM(6782) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6782)))) severity failure;
    assert RAM(6783) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6783)))) severity failure;
    assert RAM(6784) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6784)))) severity failure;
    assert RAM(6785) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6785)))) severity failure;
    assert RAM(6786) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6786)))) severity failure;
    assert RAM(6787) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6787)))) severity failure;
    assert RAM(6788) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6788)))) severity failure;
    assert RAM(6789) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6789)))) severity failure;
    assert RAM(6790) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6790)))) severity failure;
    assert RAM(6791) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6791)))) severity failure;
    assert RAM(6792) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6792)))) severity failure;
    assert RAM(6793) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6793)))) severity failure;
    assert RAM(6794) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6794)))) severity failure;
    assert RAM(6795) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6795)))) severity failure;
    assert RAM(6796) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6796)))) severity failure;
    assert RAM(6797) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6797)))) severity failure;
    assert RAM(6798) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6798)))) severity failure;
    assert RAM(6799) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6799)))) severity failure;
    assert RAM(6800) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6800)))) severity failure;
    assert RAM(6801) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6801)))) severity failure;
    assert RAM(6802) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6802)))) severity failure;
    assert RAM(6803) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6803)))) severity failure;
    assert RAM(6804) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6804)))) severity failure;
    assert RAM(6805) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6805)))) severity failure;
    assert RAM(6806) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6806)))) severity failure;
    assert RAM(6807) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6807)))) severity failure;
    assert RAM(6808) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6808)))) severity failure;
    assert RAM(6809) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6809)))) severity failure;
    assert RAM(6810) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6810)))) severity failure;
    assert RAM(6811) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6811)))) severity failure;
    assert RAM(6812) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6812)))) severity failure;
    assert RAM(6813) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6813)))) severity failure;
    assert RAM(6814) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6814)))) severity failure;
    assert RAM(6815) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6815)))) severity failure;
    assert RAM(6816) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6816)))) severity failure;
    assert RAM(6817) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6817)))) severity failure;
    assert RAM(6818) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6818)))) severity failure;
    assert RAM(6819) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6819)))) severity failure;
    assert RAM(6820) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6820)))) severity failure;
    assert RAM(6821) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6821)))) severity failure;
    assert RAM(6822) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6822)))) severity failure;
    assert RAM(6823) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6823)))) severity failure;
    assert RAM(6824) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6824)))) severity failure;
    assert RAM(6825) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6825)))) severity failure;
    assert RAM(6826) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6826)))) severity failure;
    assert RAM(6827) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6827)))) severity failure;
    assert RAM(6828) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6828)))) severity failure;
    assert RAM(6829) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6829)))) severity failure;
    assert RAM(6830) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6830)))) severity failure;
    assert RAM(6831) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6831)))) severity failure;
    assert RAM(6832) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6832)))) severity failure;
    assert RAM(6833) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6833)))) severity failure;
    assert RAM(6834) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6834)))) severity failure;
    assert RAM(6835) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6835)))) severity failure;
    assert RAM(6836) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6836)))) severity failure;
    assert RAM(6837) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6837)))) severity failure;
    assert RAM(6838) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6838)))) severity failure;
    assert RAM(6839) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6839)))) severity failure;
    assert RAM(6840) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6840)))) severity failure;
    assert RAM(6841) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6841)))) severity failure;
    assert RAM(6842) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6842)))) severity failure;
    assert RAM(6843) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6843)))) severity failure;
    assert RAM(6844) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6844)))) severity failure;
    assert RAM(6845) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6845)))) severity failure;
    assert RAM(6846) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6846)))) severity failure;
    assert RAM(6847) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6847)))) severity failure;
    assert RAM(6848) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6848)))) severity failure;
    assert RAM(6849) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6849)))) severity failure;
    assert RAM(6850) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6850)))) severity failure;
    assert RAM(6851) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6851)))) severity failure;
    assert RAM(6852) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6852)))) severity failure;
    assert RAM(6853) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6853)))) severity failure;
    assert RAM(6854) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6854)))) severity failure;
    assert RAM(6855) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6855)))) severity failure;
    assert RAM(6856) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6856)))) severity failure;
    assert RAM(6857) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6857)))) severity failure;
    assert RAM(6858) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6858)))) severity failure;
    assert RAM(6859) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6859)))) severity failure;
    assert RAM(6860) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6860)))) severity failure;
    assert RAM(6861) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6861)))) severity failure;
    assert RAM(6862) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6862)))) severity failure;
    assert RAM(6863) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6863)))) severity failure;
    assert RAM(6864) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6864)))) severity failure;
    assert RAM(6865) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6865)))) severity failure;
    assert RAM(6866) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6866)))) severity failure;
    assert RAM(6867) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6867)))) severity failure;
    assert RAM(6868) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6868)))) severity failure;
    assert RAM(6869) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6869)))) severity failure;
    assert RAM(6870) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6870)))) severity failure;
    assert RAM(6871) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6871)))) severity failure;
    assert RAM(6872) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6872)))) severity failure;
    assert RAM(6873) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6873)))) severity failure;
    assert RAM(6874) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6874)))) severity failure;
    assert RAM(6875) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6875)))) severity failure;
    assert RAM(6876) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6876)))) severity failure;
    assert RAM(6877) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6877)))) severity failure;
    assert RAM(6878) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6878)))) severity failure;
    assert RAM(6879) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6879)))) severity failure;
    assert RAM(6880) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6880)))) severity failure;
    assert RAM(6881) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6881)))) severity failure;
    assert RAM(6882) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6882)))) severity failure;
    assert RAM(6883) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6883)))) severity failure;
    assert RAM(6884) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6884)))) severity failure;
    assert RAM(6885) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6885)))) severity failure;
    assert RAM(6886) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6886)))) severity failure;
    assert RAM(6887) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6887)))) severity failure;
    assert RAM(6888) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6888)))) severity failure;
    assert RAM(6889) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6889)))) severity failure;
    assert RAM(6890) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6890)))) severity failure;
    assert RAM(6891) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6891)))) severity failure;
    assert RAM(6892) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6892)))) severity failure;
    assert RAM(6893) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6893)))) severity failure;
    assert RAM(6894) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6894)))) severity failure;
    assert RAM(6895) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6895)))) severity failure;
    assert RAM(6896) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6896)))) severity failure;
    assert RAM(6897) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6897)))) severity failure;
    assert RAM(6898) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6898)))) severity failure;
    assert RAM(6899) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6899)))) severity failure;
    assert RAM(6900) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6900)))) severity failure;
    assert RAM(6901) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6901)))) severity failure;
    assert RAM(6902) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6902)))) severity failure;
    assert RAM(6903) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6903)))) severity failure;
    assert RAM(6904) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6904)))) severity failure;
    assert RAM(6905) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6905)))) severity failure;
    assert RAM(6906) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6906)))) severity failure;
    assert RAM(6907) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6907)))) severity failure;
    assert RAM(6908) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6908)))) severity failure;
    assert RAM(6909) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6909)))) severity failure;
    assert RAM(6910) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6910)))) severity failure;
    assert RAM(6911) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6911)))) severity failure;
    assert RAM(6912) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6912)))) severity failure;
    assert RAM(6913) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6913)))) severity failure;
    assert RAM(6914) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6914)))) severity failure;
    assert RAM(6915) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6915)))) severity failure;
    assert RAM(6916) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6916)))) severity failure;
    assert RAM(6917) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6917)))) severity failure;
    assert RAM(6918) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6918)))) severity failure;
    assert RAM(6919) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6919)))) severity failure;
    assert RAM(6920) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6920)))) severity failure;
    assert RAM(6921) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6921)))) severity failure;
    assert RAM(6922) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6922)))) severity failure;
    assert RAM(6923) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6923)))) severity failure;
    assert RAM(6924) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6924)))) severity failure;
    assert RAM(6925) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6925)))) severity failure;
    assert RAM(6926) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6926)))) severity failure;
    assert RAM(6927) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6927)))) severity failure;
    assert RAM(6928) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6928)))) severity failure;
    assert RAM(6929) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6929)))) severity failure;
    assert RAM(6930) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6930)))) severity failure;
    assert RAM(6931) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6931)))) severity failure;
    assert RAM(6932) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6932)))) severity failure;
    assert RAM(6933) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6933)))) severity failure;
    assert RAM(6934) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6934)))) severity failure;
    assert RAM(6935) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6935)))) severity failure;
    assert RAM(6936) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6936)))) severity failure;
    assert RAM(6937) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6937)))) severity failure;
    assert RAM(6938) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6938)))) severity failure;
    assert RAM(6939) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6939)))) severity failure;
    assert RAM(6940) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6940)))) severity failure;
    assert RAM(6941) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6941)))) severity failure;
    assert RAM(6942) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6942)))) severity failure;
    assert RAM(6943) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6943)))) severity failure;
    assert RAM(6944) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6944)))) severity failure;
    assert RAM(6945) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6945)))) severity failure;
    assert RAM(6946) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6946)))) severity failure;
    assert RAM(6947) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6947)))) severity failure;
    assert RAM(6948) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6948)))) severity failure;
    assert RAM(6949) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6949)))) severity failure;
    assert RAM(6950) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6950)))) severity failure;
    assert RAM(6951) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6951)))) severity failure;
    assert RAM(6952) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6952)))) severity failure;
    assert RAM(6953) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6953)))) severity failure;
    assert RAM(6954) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6954)))) severity failure;
    assert RAM(6955) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6955)))) severity failure;
    assert RAM(6956) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6956)))) severity failure;
    assert RAM(6957) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6957)))) severity failure;
    assert RAM(6958) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6958)))) severity failure;
    assert RAM(6959) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6959)))) severity failure;
    assert RAM(6960) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6960)))) severity failure;
    assert RAM(6961) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6961)))) severity failure;
    assert RAM(6962) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6962)))) severity failure;
    assert RAM(6963) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6963)))) severity failure;
    assert RAM(6964) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(6964)))) severity failure;
    assert RAM(6965) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6965)))) severity failure;
    assert RAM(6966) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6966)))) severity failure;
    assert RAM(6967) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6967)))) severity failure;
    assert RAM(6968) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6968)))) severity failure;
    assert RAM(6969) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6969)))) severity failure;
    assert RAM(6970) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(6970)))) severity failure;
    assert RAM(6971) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6971)))) severity failure;
    assert RAM(6972) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6972)))) severity failure;
    assert RAM(6973) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6973)))) severity failure;
    assert RAM(6974) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6974)))) severity failure;
    assert RAM(6975) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6975)))) severity failure;
    assert RAM(6976) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6976)))) severity failure;
    assert RAM(6977) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6977)))) severity failure;
    assert RAM(6978) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6978)))) severity failure;
    assert RAM(6979) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6979)))) severity failure;
    assert RAM(6980) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(6980)))) severity failure;
    assert RAM(6981) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6981)))) severity failure;
    assert RAM(6982) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6982)))) severity failure;
    assert RAM(6983) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6983)))) severity failure;
    assert RAM(6984) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6984)))) severity failure;
    assert RAM(6985) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6985)))) severity failure;
    assert RAM(6986) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6986)))) severity failure;
    assert RAM(6987) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6987)))) severity failure;
    assert RAM(6988) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6988)))) severity failure;
    assert RAM(6989) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6989)))) severity failure;
    assert RAM(6990) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(6990)))) severity failure;
    assert RAM(6991) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6991)))) severity failure;
    assert RAM(6992) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6992)))) severity failure;
    assert RAM(6993) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6993)))) severity failure;
    assert RAM(6994) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(6994)))) severity failure;
    assert RAM(6995) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6995)))) severity failure;
    assert RAM(6996) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(6996)))) severity failure;
    assert RAM(6997) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6997)))) severity failure;
    assert RAM(6998) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6998)))) severity failure;
    assert RAM(6999) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(6999)))) severity failure;
    assert RAM(7000) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7000)))) severity failure;
    assert RAM(7001) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7001)))) severity failure;
    assert RAM(7002) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7002)))) severity failure;
    assert RAM(7003) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7003)))) severity failure;
    assert RAM(7004) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7004)))) severity failure;
    assert RAM(7005) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7005)))) severity failure;
    assert RAM(7006) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7006)))) severity failure;
    assert RAM(7007) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7007)))) severity failure;
    assert RAM(7008) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7008)))) severity failure;
    assert RAM(7009) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7009)))) severity failure;
    assert RAM(7010) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7010)))) severity failure;
    assert RAM(7011) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7011)))) severity failure;
    assert RAM(7012) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7012)))) severity failure;
    assert RAM(7013) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7013)))) severity failure;
    assert RAM(7014) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7014)))) severity failure;
    assert RAM(7015) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7015)))) severity failure;
    assert RAM(7016) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7016)))) severity failure;
    assert RAM(7017) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7017)))) severity failure;
    assert RAM(7018) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7018)))) severity failure;
    assert RAM(7019) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7019)))) severity failure;
    assert RAM(7020) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7020)))) severity failure;
    assert RAM(7021) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7021)))) severity failure;
    assert RAM(7022) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7022)))) severity failure;
    assert RAM(7023) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7023)))) severity failure;
    assert RAM(7024) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7024)))) severity failure;
    assert RAM(7025) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7025)))) severity failure;
    assert RAM(7026) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7026)))) severity failure;
    assert RAM(7027) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7027)))) severity failure;
    assert RAM(7028) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7028)))) severity failure;
    assert RAM(7029) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7029)))) severity failure;
    assert RAM(7030) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7030)))) severity failure;
    assert RAM(7031) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7031)))) severity failure;
    assert RAM(7032) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7032)))) severity failure;
    assert RAM(7033) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7033)))) severity failure;
    assert RAM(7034) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7034)))) severity failure;
    assert RAM(7035) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7035)))) severity failure;
    assert RAM(7036) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7036)))) severity failure;
    assert RAM(7037) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7037)))) severity failure;
    assert RAM(7038) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7038)))) severity failure;
    assert RAM(7039) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7039)))) severity failure;
    assert RAM(7040) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7040)))) severity failure;
    assert RAM(7041) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7041)))) severity failure;
    assert RAM(7042) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7042)))) severity failure;
    assert RAM(7043) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7043)))) severity failure;
    assert RAM(7044) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7044)))) severity failure;
    assert RAM(7045) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7045)))) severity failure;
    assert RAM(7046) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7046)))) severity failure;
    assert RAM(7047) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7047)))) severity failure;
    assert RAM(7048) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7048)))) severity failure;
    assert RAM(7049) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7049)))) severity failure;
    assert RAM(7050) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7050)))) severity failure;
    assert RAM(7051) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7051)))) severity failure;
    assert RAM(7052) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7052)))) severity failure;
    assert RAM(7053) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7053)))) severity failure;
    assert RAM(7054) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7054)))) severity failure;
    assert RAM(7055) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7055)))) severity failure;
    assert RAM(7056) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7056)))) severity failure;
    assert RAM(7057) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7057)))) severity failure;
    assert RAM(7058) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7058)))) severity failure;
    assert RAM(7059) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7059)))) severity failure;
    assert RAM(7060) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7060)))) severity failure;
    assert RAM(7061) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7061)))) severity failure;
    assert RAM(7062) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7062)))) severity failure;
    assert RAM(7063) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7063)))) severity failure;
    assert RAM(7064) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7064)))) severity failure;
    assert RAM(7065) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7065)))) severity failure;
    assert RAM(7066) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7066)))) severity failure;
    assert RAM(7067) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7067)))) severity failure;
    assert RAM(7068) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7068)))) severity failure;
    assert RAM(7069) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7069)))) severity failure;
    assert RAM(7070) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7070)))) severity failure;
    assert RAM(7071) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7071)))) severity failure;
    assert RAM(7072) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7072)))) severity failure;
    assert RAM(7073) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7073)))) severity failure;
    assert RAM(7074) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7074)))) severity failure;
    assert RAM(7075) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7075)))) severity failure;
    assert RAM(7076) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7076)))) severity failure;
    assert RAM(7077) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7077)))) severity failure;
    assert RAM(7078) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7078)))) severity failure;
    assert RAM(7079) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7079)))) severity failure;
    assert RAM(7080) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7080)))) severity failure;
    assert RAM(7081) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7081)))) severity failure;
    assert RAM(7082) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7082)))) severity failure;
    assert RAM(7083) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7083)))) severity failure;
    assert RAM(7084) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7084)))) severity failure;
    assert RAM(7085) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7085)))) severity failure;
    assert RAM(7086) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7086)))) severity failure;
    assert RAM(7087) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7087)))) severity failure;
    assert RAM(7088) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7088)))) severity failure;
    assert RAM(7089) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7089)))) severity failure;
    assert RAM(7090) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7090)))) severity failure;
    assert RAM(7091) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7091)))) severity failure;
    assert RAM(7092) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7092)))) severity failure;
    assert RAM(7093) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7093)))) severity failure;
    assert RAM(7094) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7094)))) severity failure;
    assert RAM(7095) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7095)))) severity failure;
    assert RAM(7096) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7096)))) severity failure;
    assert RAM(7097) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7097)))) severity failure;
    assert RAM(7098) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7098)))) severity failure;
    assert RAM(7099) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7099)))) severity failure;
    assert RAM(7100) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7100)))) severity failure;
    assert RAM(7101) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7101)))) severity failure;
    assert RAM(7102) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7102)))) severity failure;
    assert RAM(7103) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7103)))) severity failure;
    assert RAM(7104) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7104)))) severity failure;
    assert RAM(7105) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7105)))) severity failure;
    assert RAM(7106) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7106)))) severity failure;
    assert RAM(7107) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7107)))) severity failure;
    assert RAM(7108) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7108)))) severity failure;
    assert RAM(7109) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7109)))) severity failure;
    assert RAM(7110) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7110)))) severity failure;
    assert RAM(7111) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7111)))) severity failure;
    assert RAM(7112) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7112)))) severity failure;
    assert RAM(7113) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7113)))) severity failure;
    assert RAM(7114) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7114)))) severity failure;
    assert RAM(7115) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7115)))) severity failure;
    assert RAM(7116) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7116)))) severity failure;
    assert RAM(7117) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7117)))) severity failure;
    assert RAM(7118) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7118)))) severity failure;
    assert RAM(7119) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7119)))) severity failure;
    assert RAM(7120) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7120)))) severity failure;
    assert RAM(7121) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7121)))) severity failure;
    assert RAM(7122) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7122)))) severity failure;
    assert RAM(7123) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7123)))) severity failure;
    assert RAM(7124) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7124)))) severity failure;
    assert RAM(7125) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7125)))) severity failure;
    assert RAM(7126) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7126)))) severity failure;
    assert RAM(7127) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7127)))) severity failure;
    assert RAM(7128) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7128)))) severity failure;
    assert RAM(7129) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7129)))) severity failure;
    assert RAM(7130) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7130)))) severity failure;
    assert RAM(7131) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7131)))) severity failure;
    assert RAM(7132) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7132)))) severity failure;
    assert RAM(7133) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7133)))) severity failure;
    assert RAM(7134) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7134)))) severity failure;
    assert RAM(7135) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7135)))) severity failure;
    assert RAM(7136) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7136)))) severity failure;
    assert RAM(7137) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7137)))) severity failure;
    assert RAM(7138) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7138)))) severity failure;
    assert RAM(7139) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7139)))) severity failure;
    assert RAM(7140) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7140)))) severity failure;
    assert RAM(7141) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7141)))) severity failure;
    assert RAM(7142) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7142)))) severity failure;
    assert RAM(7143) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7143)))) severity failure;
    assert RAM(7144) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7144)))) severity failure;
    assert RAM(7145) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7145)))) severity failure;
    assert RAM(7146) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7146)))) severity failure;
    assert RAM(7147) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7147)))) severity failure;
    assert RAM(7148) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7148)))) severity failure;
    assert RAM(7149) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7149)))) severity failure;
    assert RAM(7150) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7150)))) severity failure;
    assert RAM(7151) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7151)))) severity failure;
    assert RAM(7152) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7152)))) severity failure;
    assert RAM(7153) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7153)))) severity failure;
    assert RAM(7154) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7154)))) severity failure;
    assert RAM(7155) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7155)))) severity failure;
    assert RAM(7156) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7156)))) severity failure;
    assert RAM(7157) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7157)))) severity failure;
    assert RAM(7158) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7158)))) severity failure;
    assert RAM(7159) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7159)))) severity failure;
    assert RAM(7160) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7160)))) severity failure;
    assert RAM(7161) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7161)))) severity failure;
    assert RAM(7162) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7162)))) severity failure;
    assert RAM(7163) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7163)))) severity failure;
    assert RAM(7164) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7164)))) severity failure;
    assert RAM(7165) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7165)))) severity failure;
    assert RAM(7166) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7166)))) severity failure;
    assert RAM(7167) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7167)))) severity failure;
    assert RAM(7168) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7168)))) severity failure;
    assert RAM(7169) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7169)))) severity failure;
    assert RAM(7170) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7170)))) severity failure;
    assert RAM(7171) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7171)))) severity failure;
    assert RAM(7172) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7172)))) severity failure;
    assert RAM(7173) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7173)))) severity failure;
    assert RAM(7174) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7174)))) severity failure;
    assert RAM(7175) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7175)))) severity failure;
    assert RAM(7176) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7176)))) severity failure;
    assert RAM(7177) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7177)))) severity failure;
    assert RAM(7178) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7178)))) severity failure;
    assert RAM(7179) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7179)))) severity failure;
    assert RAM(7180) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7180)))) severity failure;
    assert RAM(7181) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7181)))) severity failure;
    assert RAM(7182) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7182)))) severity failure;
    assert RAM(7183) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7183)))) severity failure;
    assert RAM(7184) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7184)))) severity failure;
    assert RAM(7185) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7185)))) severity failure;
    assert RAM(7186) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7186)))) severity failure;
    assert RAM(7187) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7187)))) severity failure;
    assert RAM(7188) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7188)))) severity failure;
    assert RAM(7189) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7189)))) severity failure;
    assert RAM(7190) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7190)))) severity failure;
    assert RAM(7191) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7191)))) severity failure;
    assert RAM(7192) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7192)))) severity failure;
    assert RAM(7193) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7193)))) severity failure;
    assert RAM(7194) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7194)))) severity failure;
    assert RAM(7195) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7195)))) severity failure;
    assert RAM(7196) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7196)))) severity failure;
    assert RAM(7197) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7197)))) severity failure;
    assert RAM(7198) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7198)))) severity failure;
    assert RAM(7199) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7199)))) severity failure;
    assert RAM(7200) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7200)))) severity failure;
    assert RAM(7201) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7201)))) severity failure;
    assert RAM(7202) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7202)))) severity failure;
    assert RAM(7203) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7203)))) severity failure;
    assert RAM(7204) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7204)))) severity failure;
    assert RAM(7205) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7205)))) severity failure;
    assert RAM(7206) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7206)))) severity failure;
    assert RAM(7207) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7207)))) severity failure;
    assert RAM(7208) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7208)))) severity failure;
    assert RAM(7209) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7209)))) severity failure;
    assert RAM(7210) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7210)))) severity failure;
    assert RAM(7211) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7211)))) severity failure;
    assert RAM(7212) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7212)))) severity failure;
    assert RAM(7213) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7213)))) severity failure;
    assert RAM(7214) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7214)))) severity failure;
    assert RAM(7215) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7215)))) severity failure;
    assert RAM(7216) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7216)))) severity failure;
    assert RAM(7217) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7217)))) severity failure;
    assert RAM(7218) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7218)))) severity failure;
    assert RAM(7219) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7219)))) severity failure;
    assert RAM(7220) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7220)))) severity failure;
    assert RAM(7221) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7221)))) severity failure;
    assert RAM(7222) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7222)))) severity failure;
    assert RAM(7223) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7223)))) severity failure;
    assert RAM(7224) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7224)))) severity failure;
    assert RAM(7225) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7225)))) severity failure;
    assert RAM(7226) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7226)))) severity failure;
    assert RAM(7227) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7227)))) severity failure;
    assert RAM(7228) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7228)))) severity failure;
    assert RAM(7229) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7229)))) severity failure;
    assert RAM(7230) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7230)))) severity failure;
    assert RAM(7231) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7231)))) severity failure;
    assert RAM(7232) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7232)))) severity failure;
    assert RAM(7233) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7233)))) severity failure;
    assert RAM(7234) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7234)))) severity failure;
    assert RAM(7235) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7235)))) severity failure;
    assert RAM(7236) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7236)))) severity failure;
    assert RAM(7237) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7237)))) severity failure;
    assert RAM(7238) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7238)))) severity failure;
    assert RAM(7239) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7239)))) severity failure;
    assert RAM(7240) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7240)))) severity failure;
    assert RAM(7241) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7241)))) severity failure;
    assert RAM(7242) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7242)))) severity failure;
    assert RAM(7243) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7243)))) severity failure;
    assert RAM(7244) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7244)))) severity failure;
    assert RAM(7245) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7245)))) severity failure;
    assert RAM(7246) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7246)))) severity failure;
    assert RAM(7247) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7247)))) severity failure;
    assert RAM(7248) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7248)))) severity failure;
    assert RAM(7249) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7249)))) severity failure;
    assert RAM(7250) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7250)))) severity failure;
    assert RAM(7251) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7251)))) severity failure;
    assert RAM(7252) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7252)))) severity failure;
    assert RAM(7253) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7253)))) severity failure;
    assert RAM(7254) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7254)))) severity failure;
    assert RAM(7255) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7255)))) severity failure;
    assert RAM(7256) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7256)))) severity failure;
    assert RAM(7257) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7257)))) severity failure;
    assert RAM(7258) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7258)))) severity failure;
    assert RAM(7259) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7259)))) severity failure;
    assert RAM(7260) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7260)))) severity failure;
    assert RAM(7261) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7261)))) severity failure;
    assert RAM(7262) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7262)))) severity failure;
    assert RAM(7263) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7263)))) severity failure;
    assert RAM(7264) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7264)))) severity failure;
    assert RAM(7265) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7265)))) severity failure;
    assert RAM(7266) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7266)))) severity failure;
    assert RAM(7267) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7267)))) severity failure;
    assert RAM(7268) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7268)))) severity failure;
    assert RAM(7269) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7269)))) severity failure;
    assert RAM(7270) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7270)))) severity failure;
    assert RAM(7271) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7271)))) severity failure;
    assert RAM(7272) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7272)))) severity failure;
    assert RAM(7273) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7273)))) severity failure;
    assert RAM(7274) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7274)))) severity failure;
    assert RAM(7275) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7275)))) severity failure;
    assert RAM(7276) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7276)))) severity failure;
    assert RAM(7277) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7277)))) severity failure;
    assert RAM(7278) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7278)))) severity failure;
    assert RAM(7279) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7279)))) severity failure;
    assert RAM(7280) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7280)))) severity failure;
    assert RAM(7281) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7281)))) severity failure;
    assert RAM(7282) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7282)))) severity failure;
    assert RAM(7283) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7283)))) severity failure;
    assert RAM(7284) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7284)))) severity failure;
    assert RAM(7285) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7285)))) severity failure;
    assert RAM(7286) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7286)))) severity failure;
    assert RAM(7287) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7287)))) severity failure;
    assert RAM(7288) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7288)))) severity failure;
    assert RAM(7289) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7289)))) severity failure;
    assert RAM(7290) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7290)))) severity failure;
    assert RAM(7291) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7291)))) severity failure;
    assert RAM(7292) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7292)))) severity failure;
    assert RAM(7293) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7293)))) severity failure;
    assert RAM(7294) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7294)))) severity failure;
    assert RAM(7295) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7295)))) severity failure;
    assert RAM(7296) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7296)))) severity failure;
    assert RAM(7297) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7297)))) severity failure;
    assert RAM(7298) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7298)))) severity failure;
    assert RAM(7299) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7299)))) severity failure;
    assert RAM(7300) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7300)))) severity failure;
    assert RAM(7301) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7301)))) severity failure;
    assert RAM(7302) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7302)))) severity failure;
    assert RAM(7303) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7303)))) severity failure;
    assert RAM(7304) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7304)))) severity failure;
    assert RAM(7305) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7305)))) severity failure;
    assert RAM(7306) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7306)))) severity failure;
    assert RAM(7307) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7307)))) severity failure;
    assert RAM(7308) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7308)))) severity failure;
    assert RAM(7309) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7309)))) severity failure;
    assert RAM(7310) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7310)))) severity failure;
    assert RAM(7311) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7311)))) severity failure;
    assert RAM(7312) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7312)))) severity failure;
    assert RAM(7313) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7313)))) severity failure;
    assert RAM(7314) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7314)))) severity failure;
    assert RAM(7315) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7315)))) severity failure;
    assert RAM(7316) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7316)))) severity failure;
    assert RAM(7317) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7317)))) severity failure;
    assert RAM(7318) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7318)))) severity failure;
    assert RAM(7319) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7319)))) severity failure;
    assert RAM(7320) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7320)))) severity failure;
    assert RAM(7321) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7321)))) severity failure;
    assert RAM(7322) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7322)))) severity failure;
    assert RAM(7323) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7323)))) severity failure;
    assert RAM(7324) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7324)))) severity failure;
    assert RAM(7325) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7325)))) severity failure;
    assert RAM(7326) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7326)))) severity failure;
    assert RAM(7327) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7327)))) severity failure;
    assert RAM(7328) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7328)))) severity failure;
    assert RAM(7329) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7329)))) severity failure;
    assert RAM(7330) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7330)))) severity failure;
    assert RAM(7331) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7331)))) severity failure;
    assert RAM(7332) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7332)))) severity failure;
    assert RAM(7333) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7333)))) severity failure;
    assert RAM(7334) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7334)))) severity failure;
    assert RAM(7335) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7335)))) severity failure;
    assert RAM(7336) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7336)))) severity failure;
    assert RAM(7337) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7337)))) severity failure;
    assert RAM(7338) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7338)))) severity failure;
    assert RAM(7339) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7339)))) severity failure;
    assert RAM(7340) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7340)))) severity failure;
    assert RAM(7341) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7341)))) severity failure;
    assert RAM(7342) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7342)))) severity failure;
    assert RAM(7343) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7343)))) severity failure;
    assert RAM(7344) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7344)))) severity failure;
    assert RAM(7345) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7345)))) severity failure;
    assert RAM(7346) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7346)))) severity failure;
    assert RAM(7347) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7347)))) severity failure;
    assert RAM(7348) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7348)))) severity failure;
    assert RAM(7349) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7349)))) severity failure;
    assert RAM(7350) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7350)))) severity failure;
    assert RAM(7351) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7351)))) severity failure;
    assert RAM(7352) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7352)))) severity failure;
    assert RAM(7353) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7353)))) severity failure;
    assert RAM(7354) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7354)))) severity failure;
    assert RAM(7355) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7355)))) severity failure;
    assert RAM(7356) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7356)))) severity failure;
    assert RAM(7357) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7357)))) severity failure;
    assert RAM(7358) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7358)))) severity failure;
    assert RAM(7359) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7359)))) severity failure;
    assert RAM(7360) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7360)))) severity failure;
    assert RAM(7361) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7361)))) severity failure;
    assert RAM(7362) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7362)))) severity failure;
    assert RAM(7363) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7363)))) severity failure;
    assert RAM(7364) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7364)))) severity failure;
    assert RAM(7365) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7365)))) severity failure;
    assert RAM(7366) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7366)))) severity failure;
    assert RAM(7367) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7367)))) severity failure;
    assert RAM(7368) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7368)))) severity failure;
    assert RAM(7369) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7369)))) severity failure;
    assert RAM(7370) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7370)))) severity failure;
    assert RAM(7371) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7371)))) severity failure;
    assert RAM(7372) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7372)))) severity failure;
    assert RAM(7373) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7373)))) severity failure;
    assert RAM(7374) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7374)))) severity failure;
    assert RAM(7375) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7375)))) severity failure;
    assert RAM(7376) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7376)))) severity failure;
    assert RAM(7377) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7377)))) severity failure;
    assert RAM(7378) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7378)))) severity failure;
    assert RAM(7379) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7379)))) severity failure;
    assert RAM(7380) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7380)))) severity failure;
    assert RAM(7381) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7381)))) severity failure;
    assert RAM(7382) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7382)))) severity failure;
    assert RAM(7383) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7383)))) severity failure;
    assert RAM(7384) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7384)))) severity failure;
    assert RAM(7385) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7385)))) severity failure;
    assert RAM(7386) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7386)))) severity failure;
    assert RAM(7387) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7387)))) severity failure;
    assert RAM(7388) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7388)))) severity failure;
    assert RAM(7389) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7389)))) severity failure;
    assert RAM(7390) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7390)))) severity failure;
    assert RAM(7391) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7391)))) severity failure;
    assert RAM(7392) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7392)))) severity failure;
    assert RAM(7393) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7393)))) severity failure;
    assert RAM(7394) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7394)))) severity failure;
    assert RAM(7395) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7395)))) severity failure;
    assert RAM(7396) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7396)))) severity failure;
    assert RAM(7397) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7397)))) severity failure;
    assert RAM(7398) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7398)))) severity failure;
    assert RAM(7399) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7399)))) severity failure;
    assert RAM(7400) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7400)))) severity failure;
    assert RAM(7401) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7401)))) severity failure;
    assert RAM(7402) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7402)))) severity failure;
    assert RAM(7403) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7403)))) severity failure;
    assert RAM(7404) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7404)))) severity failure;
    assert RAM(7405) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7405)))) severity failure;
    assert RAM(7406) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7406)))) severity failure;
    assert RAM(7407) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7407)))) severity failure;
    assert RAM(7408) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7408)))) severity failure;
    assert RAM(7409) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7409)))) severity failure;
    assert RAM(7410) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7410)))) severity failure;
    assert RAM(7411) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7411)))) severity failure;
    assert RAM(7412) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7412)))) severity failure;
    assert RAM(7413) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7413)))) severity failure;
    assert RAM(7414) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7414)))) severity failure;
    assert RAM(7415) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7415)))) severity failure;
    assert RAM(7416) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7416)))) severity failure;
    assert RAM(7417) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7417)))) severity failure;
    assert RAM(7418) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7418)))) severity failure;
    assert RAM(7419) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7419)))) severity failure;
    assert RAM(7420) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7420)))) severity failure;
    assert RAM(7421) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7421)))) severity failure;
    assert RAM(7422) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7422)))) severity failure;
    assert RAM(7423) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7423)))) severity failure;
    assert RAM(7424) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7424)))) severity failure;
    assert RAM(7425) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7425)))) severity failure;
    assert RAM(7426) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7426)))) severity failure;
    assert RAM(7427) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7427)))) severity failure;
    assert RAM(7428) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7428)))) severity failure;
    assert RAM(7429) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7429)))) severity failure;
    assert RAM(7430) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7430)))) severity failure;
    assert RAM(7431) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7431)))) severity failure;
    assert RAM(7432) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7432)))) severity failure;
    assert RAM(7433) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7433)))) severity failure;
    assert RAM(7434) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7434)))) severity failure;
    assert RAM(7435) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7435)))) severity failure;
    assert RAM(7436) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7436)))) severity failure;
    assert RAM(7437) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7437)))) severity failure;
    assert RAM(7438) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7438)))) severity failure;
    assert RAM(7439) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7439)))) severity failure;
    assert RAM(7440) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7440)))) severity failure;
    assert RAM(7441) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7441)))) severity failure;
    assert RAM(7442) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7442)))) severity failure;
    assert RAM(7443) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7443)))) severity failure;
    assert RAM(7444) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7444)))) severity failure;
    assert RAM(7445) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7445)))) severity failure;
    assert RAM(7446) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7446)))) severity failure;
    assert RAM(7447) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7447)))) severity failure;
    assert RAM(7448) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7448)))) severity failure;
    assert RAM(7449) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7449)))) severity failure;
    assert RAM(7450) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7450)))) severity failure;
    assert RAM(7451) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7451)))) severity failure;
    assert RAM(7452) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7452)))) severity failure;
    assert RAM(7453) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7453)))) severity failure;
    assert RAM(7454) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7454)))) severity failure;
    assert RAM(7455) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7455)))) severity failure;
    assert RAM(7456) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7456)))) severity failure;
    assert RAM(7457) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7457)))) severity failure;
    assert RAM(7458) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7458)))) severity failure;
    assert RAM(7459) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7459)))) severity failure;
    assert RAM(7460) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7460)))) severity failure;
    assert RAM(7461) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7461)))) severity failure;
    assert RAM(7462) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7462)))) severity failure;
    assert RAM(7463) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7463)))) severity failure;
    assert RAM(7464) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7464)))) severity failure;
    assert RAM(7465) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7465)))) severity failure;
    assert RAM(7466) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7466)))) severity failure;
    assert RAM(7467) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7467)))) severity failure;
    assert RAM(7468) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7468)))) severity failure;
    assert RAM(7469) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7469)))) severity failure;
    assert RAM(7470) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7470)))) severity failure;
    assert RAM(7471) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7471)))) severity failure;
    assert RAM(7472) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7472)))) severity failure;
    assert RAM(7473) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7473)))) severity failure;
    assert RAM(7474) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7474)))) severity failure;
    assert RAM(7475) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7475)))) severity failure;
    assert RAM(7476) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7476)))) severity failure;
    assert RAM(7477) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7477)))) severity failure;
    assert RAM(7478) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7478)))) severity failure;
    assert RAM(7479) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7479)))) severity failure;
    assert RAM(7480) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7480)))) severity failure;
    assert RAM(7481) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7481)))) severity failure;
    assert RAM(7482) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7482)))) severity failure;
    assert RAM(7483) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7483)))) severity failure;
    assert RAM(7484) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7484)))) severity failure;
    assert RAM(7485) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7485)))) severity failure;
    assert RAM(7486) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7486)))) severity failure;
    assert RAM(7487) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7487)))) severity failure;
    assert RAM(7488) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7488)))) severity failure;
    assert RAM(7489) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7489)))) severity failure;
    assert RAM(7490) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7490)))) severity failure;
    assert RAM(7491) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7491)))) severity failure;
    assert RAM(7492) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7492)))) severity failure;
    assert RAM(7493) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7493)))) severity failure;
    assert RAM(7494) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7494)))) severity failure;
    assert RAM(7495) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7495)))) severity failure;
    assert RAM(7496) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7496)))) severity failure;
    assert RAM(7497) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7497)))) severity failure;
    assert RAM(7498) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7498)))) severity failure;
    assert RAM(7499) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7499)))) severity failure;
    assert RAM(7500) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7500)))) severity failure;
    assert RAM(7501) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7501)))) severity failure;
    assert RAM(7502) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7502)))) severity failure;
    assert RAM(7503) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7503)))) severity failure;
    assert RAM(7504) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7504)))) severity failure;
    assert RAM(7505) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7505)))) severity failure;
    assert RAM(7506) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7506)))) severity failure;
    assert RAM(7507) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7507)))) severity failure;
    assert RAM(7508) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7508)))) severity failure;
    assert RAM(7509) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7509)))) severity failure;
    assert RAM(7510) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7510)))) severity failure;
    assert RAM(7511) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7511)))) severity failure;
    assert RAM(7512) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7512)))) severity failure;
    assert RAM(7513) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7513)))) severity failure;
    assert RAM(7514) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7514)))) severity failure;
    assert RAM(7515) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7515)))) severity failure;
    assert RAM(7516) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7516)))) severity failure;
    assert RAM(7517) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7517)))) severity failure;
    assert RAM(7518) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7518)))) severity failure;
    assert RAM(7519) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7519)))) severity failure;
    assert RAM(7520) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7520)))) severity failure;
    assert RAM(7521) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7521)))) severity failure;
    assert RAM(7522) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7522)))) severity failure;
    assert RAM(7523) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7523)))) severity failure;
    assert RAM(7524) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7524)))) severity failure;
    assert RAM(7525) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7525)))) severity failure;
    assert RAM(7526) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7526)))) severity failure;
    assert RAM(7527) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7527)))) severity failure;
    assert RAM(7528) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7528)))) severity failure;
    assert RAM(7529) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7529)))) severity failure;
    assert RAM(7530) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7530)))) severity failure;
    assert RAM(7531) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7531)))) severity failure;
    assert RAM(7532) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7532)))) severity failure;
    assert RAM(7533) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7533)))) severity failure;
    assert RAM(7534) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7534)))) severity failure;
    assert RAM(7535) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7535)))) severity failure;
    assert RAM(7536) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7536)))) severity failure;
    assert RAM(7537) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7537)))) severity failure;
    assert RAM(7538) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7538)))) severity failure;
    assert RAM(7539) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7539)))) severity failure;
    assert RAM(7540) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7540)))) severity failure;
    assert RAM(7541) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7541)))) severity failure;
    assert RAM(7542) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7542)))) severity failure;
    assert RAM(7543) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7543)))) severity failure;
    assert RAM(7544) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7544)))) severity failure;
    assert RAM(7545) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7545)))) severity failure;
    assert RAM(7546) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7546)))) severity failure;
    assert RAM(7547) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7547)))) severity failure;
    assert RAM(7548) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7548)))) severity failure;
    assert RAM(7549) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7549)))) severity failure;
    assert RAM(7550) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7550)))) severity failure;
    assert RAM(7551) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7551)))) severity failure;
    assert RAM(7552) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7552)))) severity failure;
    assert RAM(7553) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7553)))) severity failure;
    assert RAM(7554) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7554)))) severity failure;
    assert RAM(7555) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7555)))) severity failure;
    assert RAM(7556) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7556)))) severity failure;
    assert RAM(7557) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7557)))) severity failure;
    assert RAM(7558) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7558)))) severity failure;
    assert RAM(7559) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7559)))) severity failure;
    assert RAM(7560) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7560)))) severity failure;
    assert RAM(7561) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7561)))) severity failure;
    assert RAM(7562) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7562)))) severity failure;
    assert RAM(7563) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7563)))) severity failure;
    assert RAM(7564) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7564)))) severity failure;
    assert RAM(7565) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7565)))) severity failure;
    assert RAM(7566) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7566)))) severity failure;
    assert RAM(7567) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7567)))) severity failure;
    assert RAM(7568) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7568)))) severity failure;
    assert RAM(7569) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7569)))) severity failure;
    assert RAM(7570) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7570)))) severity failure;
    assert RAM(7571) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7571)))) severity failure;
    assert RAM(7572) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7572)))) severity failure;
    assert RAM(7573) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7573)))) severity failure;
    assert RAM(7574) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7574)))) severity failure;
    assert RAM(7575) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7575)))) severity failure;
    assert RAM(7576) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7576)))) severity failure;
    assert RAM(7577) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7577)))) severity failure;
    assert RAM(7578) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7578)))) severity failure;
    assert RAM(7579) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7579)))) severity failure;
    assert RAM(7580) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7580)))) severity failure;
    assert RAM(7581) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7581)))) severity failure;
    assert RAM(7582) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7582)))) severity failure;
    assert RAM(7583) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7583)))) severity failure;
    assert RAM(7584) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7584)))) severity failure;
    assert RAM(7585) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7585)))) severity failure;
    assert RAM(7586) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7586)))) severity failure;
    assert RAM(7587) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7587)))) severity failure;
    assert RAM(7588) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7588)))) severity failure;
    assert RAM(7589) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7589)))) severity failure;
    assert RAM(7590) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7590)))) severity failure;
    assert RAM(7591) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7591)))) severity failure;
    assert RAM(7592) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7592)))) severity failure;
    assert RAM(7593) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7593)))) severity failure;
    assert RAM(7594) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7594)))) severity failure;
    assert RAM(7595) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7595)))) severity failure;
    assert RAM(7596) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7596)))) severity failure;
    assert RAM(7597) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7597)))) severity failure;
    assert RAM(7598) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7598)))) severity failure;
    assert RAM(7599) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7599)))) severity failure;
    assert RAM(7600) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7600)))) severity failure;
    assert RAM(7601) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7601)))) severity failure;
    assert RAM(7602) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7602)))) severity failure;
    assert RAM(7603) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7603)))) severity failure;
    assert RAM(7604) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7604)))) severity failure;
    assert RAM(7605) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7605)))) severity failure;
    assert RAM(7606) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7606)))) severity failure;
    assert RAM(7607) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7607)))) severity failure;
    assert RAM(7608) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7608)))) severity failure;
    assert RAM(7609) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7609)))) severity failure;
    assert RAM(7610) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7610)))) severity failure;
    assert RAM(7611) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7611)))) severity failure;
    assert RAM(7612) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7612)))) severity failure;
    assert RAM(7613) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7613)))) severity failure;
    assert RAM(7614) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7614)))) severity failure;
    assert RAM(7615) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7615)))) severity failure;
    assert RAM(7616) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7616)))) severity failure;
    assert RAM(7617) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7617)))) severity failure;
    assert RAM(7618) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7618)))) severity failure;
    assert RAM(7619) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7619)))) severity failure;
    assert RAM(7620) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7620)))) severity failure;
    assert RAM(7621) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7621)))) severity failure;
    assert RAM(7622) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7622)))) severity failure;
    assert RAM(7623) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7623)))) severity failure;
    assert RAM(7624) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7624)))) severity failure;
    assert RAM(7625) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7625)))) severity failure;
    assert RAM(7626) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7626)))) severity failure;
    assert RAM(7627) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7627)))) severity failure;
    assert RAM(7628) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7628)))) severity failure;
    assert RAM(7629) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7629)))) severity failure;
    assert RAM(7630) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7630)))) severity failure;
    assert RAM(7631) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7631)))) severity failure;
    assert RAM(7632) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7632)))) severity failure;
    assert RAM(7633) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7633)))) severity failure;
    assert RAM(7634) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7634)))) severity failure;
    assert RAM(7635) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7635)))) severity failure;
    assert RAM(7636) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7636)))) severity failure;
    assert RAM(7637) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7637)))) severity failure;
    assert RAM(7638) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7638)))) severity failure;
    assert RAM(7639) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7639)))) severity failure;
    assert RAM(7640) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7640)))) severity failure;
    assert RAM(7641) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7641)))) severity failure;
    assert RAM(7642) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7642)))) severity failure;
    assert RAM(7643) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7643)))) severity failure;
    assert RAM(7644) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7644)))) severity failure;
    assert RAM(7645) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7645)))) severity failure;
    assert RAM(7646) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7646)))) severity failure;
    assert RAM(7647) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7647)))) severity failure;
    assert RAM(7648) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7648)))) severity failure;
    assert RAM(7649) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7649)))) severity failure;
    assert RAM(7650) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7650)))) severity failure;
    assert RAM(7651) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7651)))) severity failure;
    assert RAM(7652) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7652)))) severity failure;
    assert RAM(7653) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7653)))) severity failure;
    assert RAM(7654) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7654)))) severity failure;
    assert RAM(7655) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7655)))) severity failure;
    assert RAM(7656) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7656)))) severity failure;
    assert RAM(7657) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7657)))) severity failure;
    assert RAM(7658) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7658)))) severity failure;
    assert RAM(7659) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7659)))) severity failure;
    assert RAM(7660) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7660)))) severity failure;
    assert RAM(7661) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7661)))) severity failure;
    assert RAM(7662) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7662)))) severity failure;
    assert RAM(7663) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7663)))) severity failure;
    assert RAM(7664) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7664)))) severity failure;
    assert RAM(7665) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7665)))) severity failure;
    assert RAM(7666) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7666)))) severity failure;
    assert RAM(7667) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7667)))) severity failure;
    assert RAM(7668) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7668)))) severity failure;
    assert RAM(7669) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7669)))) severity failure;
    assert RAM(7670) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7670)))) severity failure;
    assert RAM(7671) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7671)))) severity failure;
    assert RAM(7672) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7672)))) severity failure;
    assert RAM(7673) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7673)))) severity failure;
    assert RAM(7674) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7674)))) severity failure;
    assert RAM(7675) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7675)))) severity failure;
    assert RAM(7676) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7676)))) severity failure;
    assert RAM(7677) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7677)))) severity failure;
    assert RAM(7678) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7678)))) severity failure;
    assert RAM(7679) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7679)))) severity failure;
    assert RAM(7680) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7680)))) severity failure;
    assert RAM(7681) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7681)))) severity failure;
    assert RAM(7682) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7682)))) severity failure;
    assert RAM(7683) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7683)))) severity failure;
    assert RAM(7684) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7684)))) severity failure;
    assert RAM(7685) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7685)))) severity failure;
    assert RAM(7686) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7686)))) severity failure;
    assert RAM(7687) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7687)))) severity failure;
    assert RAM(7688) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7688)))) severity failure;
    assert RAM(7689) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7689)))) severity failure;
    assert RAM(7690) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7690)))) severity failure;
    assert RAM(7691) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7691)))) severity failure;
    assert RAM(7692) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7692)))) severity failure;
    assert RAM(7693) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7693)))) severity failure;
    assert RAM(7694) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7694)))) severity failure;
    assert RAM(7695) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7695)))) severity failure;
    assert RAM(7696) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7696)))) severity failure;
    assert RAM(7697) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7697)))) severity failure;
    assert RAM(7698) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7698)))) severity failure;
    assert RAM(7699) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7699)))) severity failure;
    assert RAM(7700) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7700)))) severity failure;
    assert RAM(7701) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7701)))) severity failure;
    assert RAM(7702) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7702)))) severity failure;
    assert RAM(7703) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7703)))) severity failure;
    assert RAM(7704) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7704)))) severity failure;
    assert RAM(7705) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7705)))) severity failure;
    assert RAM(7706) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7706)))) severity failure;
    assert RAM(7707) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7707)))) severity failure;
    assert RAM(7708) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7708)))) severity failure;
    assert RAM(7709) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7709)))) severity failure;
    assert RAM(7710) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7710)))) severity failure;
    assert RAM(7711) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7711)))) severity failure;
    assert RAM(7712) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7712)))) severity failure;
    assert RAM(7713) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7713)))) severity failure;
    assert RAM(7714) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7714)))) severity failure;
    assert RAM(7715) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7715)))) severity failure;
    assert RAM(7716) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7716)))) severity failure;
    assert RAM(7717) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7717)))) severity failure;
    assert RAM(7718) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7718)))) severity failure;
    assert RAM(7719) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7719)))) severity failure;
    assert RAM(7720) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7720)))) severity failure;
    assert RAM(7721) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7721)))) severity failure;
    assert RAM(7722) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7722)))) severity failure;
    assert RAM(7723) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7723)))) severity failure;
    assert RAM(7724) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7724)))) severity failure;
    assert RAM(7725) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7725)))) severity failure;
    assert RAM(7726) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7726)))) severity failure;
    assert RAM(7727) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7727)))) severity failure;
    assert RAM(7728) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7728)))) severity failure;
    assert RAM(7729) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7729)))) severity failure;
    assert RAM(7730) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7730)))) severity failure;
    assert RAM(7731) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7731)))) severity failure;
    assert RAM(7732) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7732)))) severity failure;
    assert RAM(7733) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7733)))) severity failure;
    assert RAM(7734) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7734)))) severity failure;
    assert RAM(7735) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7735)))) severity failure;
    assert RAM(7736) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7736)))) severity failure;
    assert RAM(7737) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7737)))) severity failure;
    assert RAM(7738) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7738)))) severity failure;
    assert RAM(7739) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7739)))) severity failure;
    assert RAM(7740) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7740)))) severity failure;
    assert RAM(7741) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7741)))) severity failure;
    assert RAM(7742) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7742)))) severity failure;
    assert RAM(7743) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7743)))) severity failure;
    assert RAM(7744) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7744)))) severity failure;
    assert RAM(7745) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7745)))) severity failure;
    assert RAM(7746) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7746)))) severity failure;
    assert RAM(7747) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7747)))) severity failure;
    assert RAM(7748) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7748)))) severity failure;
    assert RAM(7749) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7749)))) severity failure;
    assert RAM(7750) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7750)))) severity failure;
    assert RAM(7751) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7751)))) severity failure;
    assert RAM(7752) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7752)))) severity failure;
    assert RAM(7753) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7753)))) severity failure;
    assert RAM(7754) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7754)))) severity failure;
    assert RAM(7755) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7755)))) severity failure;
    assert RAM(7756) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7756)))) severity failure;
    assert RAM(7757) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7757)))) severity failure;
    assert RAM(7758) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7758)))) severity failure;
    assert RAM(7759) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7759)))) severity failure;
    assert RAM(7760) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7760)))) severity failure;
    assert RAM(7761) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7761)))) severity failure;
    assert RAM(7762) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7762)))) severity failure;
    assert RAM(7763) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7763)))) severity failure;
    assert RAM(7764) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7764)))) severity failure;
    assert RAM(7765) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7765)))) severity failure;
    assert RAM(7766) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7766)))) severity failure;
    assert RAM(7767) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7767)))) severity failure;
    assert RAM(7768) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7768)))) severity failure;
    assert RAM(7769) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7769)))) severity failure;
    assert RAM(7770) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7770)))) severity failure;
    assert RAM(7771) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7771)))) severity failure;
    assert RAM(7772) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7772)))) severity failure;
    assert RAM(7773) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7773)))) severity failure;
    assert RAM(7774) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7774)))) severity failure;
    assert RAM(7775) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7775)))) severity failure;
    assert RAM(7776) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7776)))) severity failure;
    assert RAM(7777) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7777)))) severity failure;
    assert RAM(7778) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7778)))) severity failure;
    assert RAM(7779) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7779)))) severity failure;
    assert RAM(7780) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7780)))) severity failure;
    assert RAM(7781) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7781)))) severity failure;
    assert RAM(7782) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7782)))) severity failure;
    assert RAM(7783) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7783)))) severity failure;
    assert RAM(7784) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7784)))) severity failure;
    assert RAM(7785) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7785)))) severity failure;
    assert RAM(7786) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7786)))) severity failure;
    assert RAM(7787) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7787)))) severity failure;
    assert RAM(7788) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7788)))) severity failure;
    assert RAM(7789) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7789)))) severity failure;
    assert RAM(7790) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7790)))) severity failure;
    assert RAM(7791) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7791)))) severity failure;
    assert RAM(7792) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7792)))) severity failure;
    assert RAM(7793) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7793)))) severity failure;
    assert RAM(7794) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7794)))) severity failure;
    assert RAM(7795) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7795)))) severity failure;
    assert RAM(7796) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7796)))) severity failure;
    assert RAM(7797) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7797)))) severity failure;
    assert RAM(7798) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7798)))) severity failure;
    assert RAM(7799) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7799)))) severity failure;
    assert RAM(7800) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7800)))) severity failure;
    assert RAM(7801) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7801)))) severity failure;
    assert RAM(7802) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7802)))) severity failure;
    assert RAM(7803) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7803)))) severity failure;
    assert RAM(7804) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7804)))) severity failure;
    assert RAM(7805) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7805)))) severity failure;
    assert RAM(7806) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7806)))) severity failure;
    assert RAM(7807) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7807)))) severity failure;
    assert RAM(7808) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7808)))) severity failure;
    assert RAM(7809) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7809)))) severity failure;
    assert RAM(7810) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7810)))) severity failure;
    assert RAM(7811) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7811)))) severity failure;
    assert RAM(7812) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7812)))) severity failure;
    assert RAM(7813) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7813)))) severity failure;
    assert RAM(7814) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7814)))) severity failure;
    assert RAM(7815) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7815)))) severity failure;
    assert RAM(7816) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7816)))) severity failure;
    assert RAM(7817) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7817)))) severity failure;
    assert RAM(7818) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7818)))) severity failure;
    assert RAM(7819) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7819)))) severity failure;
    assert RAM(7820) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7820)))) severity failure;
    assert RAM(7821) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7821)))) severity failure;
    assert RAM(7822) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7822)))) severity failure;
    assert RAM(7823) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7823)))) severity failure;
    assert RAM(7824) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7824)))) severity failure;
    assert RAM(7825) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7825)))) severity failure;
    assert RAM(7826) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7826)))) severity failure;
    assert RAM(7827) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7827)))) severity failure;
    assert RAM(7828) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7828)))) severity failure;
    assert RAM(7829) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7829)))) severity failure;
    assert RAM(7830) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7830)))) severity failure;
    assert RAM(7831) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7831)))) severity failure;
    assert RAM(7832) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7832)))) severity failure;
    assert RAM(7833) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7833)))) severity failure;
    assert RAM(7834) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7834)))) severity failure;
    assert RAM(7835) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7835)))) severity failure;
    assert RAM(7836) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7836)))) severity failure;
    assert RAM(7837) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7837)))) severity failure;
    assert RAM(7838) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7838)))) severity failure;
    assert RAM(7839) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7839)))) severity failure;
    assert RAM(7840) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7840)))) severity failure;
    assert RAM(7841) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7841)))) severity failure;
    assert RAM(7842) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7842)))) severity failure;
    assert RAM(7843) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7843)))) severity failure;
    assert RAM(7844) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7844)))) severity failure;
    assert RAM(7845) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7845)))) severity failure;
    assert RAM(7846) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7846)))) severity failure;
    assert RAM(7847) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7847)))) severity failure;
    assert RAM(7848) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7848)))) severity failure;
    assert RAM(7849) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7849)))) severity failure;
    assert RAM(7850) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7850)))) severity failure;
    assert RAM(7851) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7851)))) severity failure;
    assert RAM(7852) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7852)))) severity failure;
    assert RAM(7853) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7853)))) severity failure;
    assert RAM(7854) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7854)))) severity failure;
    assert RAM(7855) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7855)))) severity failure;
    assert RAM(7856) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7856)))) severity failure;
    assert RAM(7857) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7857)))) severity failure;
    assert RAM(7858) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7858)))) severity failure;
    assert RAM(7859) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7859)))) severity failure;
    assert RAM(7860) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7860)))) severity failure;
    assert RAM(7861) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7861)))) severity failure;
    assert RAM(7862) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7862)))) severity failure;
    assert RAM(7863) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7863)))) severity failure;
    assert RAM(7864) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7864)))) severity failure;
    assert RAM(7865) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7865)))) severity failure;
    assert RAM(7866) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7866)))) severity failure;
    assert RAM(7867) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7867)))) severity failure;
    assert RAM(7868) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7868)))) severity failure;
    assert RAM(7869) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7869)))) severity failure;
    assert RAM(7870) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7870)))) severity failure;
    assert RAM(7871) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7871)))) severity failure;
    assert RAM(7872) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7872)))) severity failure;
    assert RAM(7873) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7873)))) severity failure;
    assert RAM(7874) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7874)))) severity failure;
    assert RAM(7875) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7875)))) severity failure;
    assert RAM(7876) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7876)))) severity failure;
    assert RAM(7877) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7877)))) severity failure;
    assert RAM(7878) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7878)))) severity failure;
    assert RAM(7879) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7879)))) severity failure;
    assert RAM(7880) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7880)))) severity failure;
    assert RAM(7881) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7881)))) severity failure;
    assert RAM(7882) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7882)))) severity failure;
    assert RAM(7883) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7883)))) severity failure;
    assert RAM(7884) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7884)))) severity failure;
    assert RAM(7885) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7885)))) severity failure;
    assert RAM(7886) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7886)))) severity failure;
    assert RAM(7887) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7887)))) severity failure;
    assert RAM(7888) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7888)))) severity failure;
    assert RAM(7889) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7889)))) severity failure;
    assert RAM(7890) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7890)))) severity failure;
    assert RAM(7891) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7891)))) severity failure;
    assert RAM(7892) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7892)))) severity failure;
    assert RAM(7893) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7893)))) severity failure;
    assert RAM(7894) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7894)))) severity failure;
    assert RAM(7895) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7895)))) severity failure;
    assert RAM(7896) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7896)))) severity failure;
    assert RAM(7897) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7897)))) severity failure;
    assert RAM(7898) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7898)))) severity failure;
    assert RAM(7899) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7899)))) severity failure;
    assert RAM(7900) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7900)))) severity failure;
    assert RAM(7901) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7901)))) severity failure;
    assert RAM(7902) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7902)))) severity failure;
    assert RAM(7903) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7903)))) severity failure;
    assert RAM(7904) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7904)))) severity failure;
    assert RAM(7905) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7905)))) severity failure;
    assert RAM(7906) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7906)))) severity failure;
    assert RAM(7907) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7907)))) severity failure;
    assert RAM(7908) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7908)))) severity failure;
    assert RAM(7909) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7909)))) severity failure;
    assert RAM(7910) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7910)))) severity failure;
    assert RAM(7911) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7911)))) severity failure;
    assert RAM(7912) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7912)))) severity failure;
    assert RAM(7913) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7913)))) severity failure;
    assert RAM(7914) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7914)))) severity failure;
    assert RAM(7915) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7915)))) severity failure;
    assert RAM(7916) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7916)))) severity failure;
    assert RAM(7917) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7917)))) severity failure;
    assert RAM(7918) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7918)))) severity failure;
    assert RAM(7919) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7919)))) severity failure;
    assert RAM(7920) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7920)))) severity failure;
    assert RAM(7921) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7921)))) severity failure;
    assert RAM(7922) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7922)))) severity failure;
    assert RAM(7923) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7923)))) severity failure;
    assert RAM(7924) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7924)))) severity failure;
    assert RAM(7925) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7925)))) severity failure;
    assert RAM(7926) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7926)))) severity failure;
    assert RAM(7927) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7927)))) severity failure;
    assert RAM(7928) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7928)))) severity failure;
    assert RAM(7929) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7929)))) severity failure;
    assert RAM(7930) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7930)))) severity failure;
    assert RAM(7931) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7931)))) severity failure;
    assert RAM(7932) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7932)))) severity failure;
    assert RAM(7933) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7933)))) severity failure;
    assert RAM(7934) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7934)))) severity failure;
    assert RAM(7935) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7935)))) severity failure;
    assert RAM(7936) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7936)))) severity failure;
    assert RAM(7937) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7937)))) severity failure;
    assert RAM(7938) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7938)))) severity failure;
    assert RAM(7939) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7939)))) severity failure;
    assert RAM(7940) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7940)))) severity failure;
    assert RAM(7941) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7941)))) severity failure;
    assert RAM(7942) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7942)))) severity failure;
    assert RAM(7943) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7943)))) severity failure;
    assert RAM(7944) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7944)))) severity failure;
    assert RAM(7945) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7945)))) severity failure;
    assert RAM(7946) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7946)))) severity failure;
    assert RAM(7947) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7947)))) severity failure;
    assert RAM(7948) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7948)))) severity failure;
    assert RAM(7949) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7949)))) severity failure;
    assert RAM(7950) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7950)))) severity failure;
    assert RAM(7951) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7951)))) severity failure;
    assert RAM(7952) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7952)))) severity failure;
    assert RAM(7953) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7953)))) severity failure;
    assert RAM(7954) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7954)))) severity failure;
    assert RAM(7955) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7955)))) severity failure;
    assert RAM(7956) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7956)))) severity failure;
    assert RAM(7957) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7957)))) severity failure;
    assert RAM(7958) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7958)))) severity failure;
    assert RAM(7959) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7959)))) severity failure;
    assert RAM(7960) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7960)))) severity failure;
    assert RAM(7961) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7961)))) severity failure;
    assert RAM(7962) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7962)))) severity failure;
    assert RAM(7963) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(7963)))) severity failure;
    assert RAM(7964) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7964)))) severity failure;
    assert RAM(7965) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7965)))) severity failure;
    assert RAM(7966) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7966)))) severity failure;
    assert RAM(7967) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7967)))) severity failure;
    assert RAM(7968) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7968)))) severity failure;
    assert RAM(7969) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7969)))) severity failure;
    assert RAM(7970) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(7970)))) severity failure;
    assert RAM(7971) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7971)))) severity failure;
    assert RAM(7972) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7972)))) severity failure;
    assert RAM(7973) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7973)))) severity failure;
    assert RAM(7974) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7974)))) severity failure;
    assert RAM(7975) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7975)))) severity failure;
    assert RAM(7976) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7976)))) severity failure;
    assert RAM(7977) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7977)))) severity failure;
    assert RAM(7978) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7978)))) severity failure;
    assert RAM(7979) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7979)))) severity failure;
    assert RAM(7980) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7980)))) severity failure;
    assert RAM(7981) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7981)))) severity failure;
    assert RAM(7982) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7982)))) severity failure;
    assert RAM(7983) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7983)))) severity failure;
    assert RAM(7984) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7984)))) severity failure;
    assert RAM(7985) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7985)))) severity failure;
    assert RAM(7986) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7986)))) severity failure;
    assert RAM(7987) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7987)))) severity failure;
    assert RAM(7988) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7988)))) severity failure;
    assert RAM(7989) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7989)))) severity failure;
    assert RAM(7990) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(7990)))) severity failure;
    assert RAM(7991) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7991)))) severity failure;
    assert RAM(7992) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7992)))) severity failure;
    assert RAM(7993) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7993)))) severity failure;
    assert RAM(7994) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7994)))) severity failure;
    assert RAM(7995) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7995)))) severity failure;
    assert RAM(7996) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(7996)))) severity failure;
    assert RAM(7997) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(7997)))) severity failure;
    assert RAM(7998) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(7998)))) severity failure;
    assert RAM(7999) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(7999)))) severity failure;
    assert RAM(8000) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8000)))) severity failure;
    assert RAM(8001) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8001)))) severity failure;
    assert RAM(8002) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8002)))) severity failure;
    assert RAM(8003) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8003)))) severity failure;
    assert RAM(8004) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8004)))) severity failure;
    assert RAM(8005) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8005)))) severity failure;
    assert RAM(8006) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8006)))) severity failure;
    assert RAM(8007) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8007)))) severity failure;
    assert RAM(8008) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8008)))) severity failure;
    assert RAM(8009) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8009)))) severity failure;
    assert RAM(8010) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8010)))) severity failure;
    assert RAM(8011) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8011)))) severity failure;
    assert RAM(8012) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8012)))) severity failure;
    assert RAM(8013) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8013)))) severity failure;
    assert RAM(8014) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8014)))) severity failure;
    assert RAM(8015) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8015)))) severity failure;
    assert RAM(8016) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8016)))) severity failure;
    assert RAM(8017) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8017)))) severity failure;
    assert RAM(8018) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8018)))) severity failure;
    assert RAM(8019) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8019)))) severity failure;
    assert RAM(8020) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8020)))) severity failure;
    assert RAM(8021) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8021)))) severity failure;
    assert RAM(8022) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8022)))) severity failure;
    assert RAM(8023) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8023)))) severity failure;
    assert RAM(8024) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8024)))) severity failure;
    assert RAM(8025) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8025)))) severity failure;
    assert RAM(8026) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8026)))) severity failure;
    assert RAM(8027) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8027)))) severity failure;
    assert RAM(8028) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8028)))) severity failure;
    assert RAM(8029) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8029)))) severity failure;
    assert RAM(8030) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8030)))) severity failure;
    assert RAM(8031) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8031)))) severity failure;
    assert RAM(8032) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8032)))) severity failure;
    assert RAM(8033) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8033)))) severity failure;
    assert RAM(8034) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8034)))) severity failure;
    assert RAM(8035) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8035)))) severity failure;
    assert RAM(8036) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8036)))) severity failure;
    assert RAM(8037) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8037)))) severity failure;
    assert RAM(8038) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8038)))) severity failure;
    assert RAM(8039) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8039)))) severity failure;
    assert RAM(8040) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8040)))) severity failure;
    assert RAM(8041) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8041)))) severity failure;
    assert RAM(8042) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8042)))) severity failure;
    assert RAM(8043) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8043)))) severity failure;
    assert RAM(8044) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8044)))) severity failure;
    assert RAM(8045) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8045)))) severity failure;
    assert RAM(8046) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8046)))) severity failure;
    assert RAM(8047) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8047)))) severity failure;
    assert RAM(8048) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8048)))) severity failure;
    assert RAM(8049) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8049)))) severity failure;
    assert RAM(8050) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8050)))) severity failure;
    assert RAM(8051) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8051)))) severity failure;
    assert RAM(8052) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8052)))) severity failure;
    assert RAM(8053) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8053)))) severity failure;
    assert RAM(8054) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8054)))) severity failure;
    assert RAM(8055) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8055)))) severity failure;
    assert RAM(8056) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8056)))) severity failure;
    assert RAM(8057) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8057)))) severity failure;
    assert RAM(8058) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8058)))) severity failure;
    assert RAM(8059) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8059)))) severity failure;
    assert RAM(8060) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8060)))) severity failure;
    assert RAM(8061) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8061)))) severity failure;
    assert RAM(8062) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8062)))) severity failure;
    assert RAM(8063) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8063)))) severity failure;
    assert RAM(8064) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8064)))) severity failure;
    assert RAM(8065) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8065)))) severity failure;
    assert RAM(8066) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8066)))) severity failure;
    assert RAM(8067) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8067)))) severity failure;
    assert RAM(8068) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8068)))) severity failure;
    assert RAM(8069) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8069)))) severity failure;
    assert RAM(8070) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8070)))) severity failure;
    assert RAM(8071) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8071)))) severity failure;
    assert RAM(8072) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8072)))) severity failure;
    assert RAM(8073) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8073)))) severity failure;
    assert RAM(8074) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8074)))) severity failure;
    assert RAM(8075) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8075)))) severity failure;
    assert RAM(8076) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8076)))) severity failure;
    assert RAM(8077) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8077)))) severity failure;
    assert RAM(8078) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8078)))) severity failure;
    assert RAM(8079) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8079)))) severity failure;
    assert RAM(8080) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8080)))) severity failure;
    assert RAM(8081) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8081)))) severity failure;
    assert RAM(8082) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8082)))) severity failure;
    assert RAM(8083) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8083)))) severity failure;
    assert RAM(8084) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8084)))) severity failure;
    assert RAM(8085) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8085)))) severity failure;
    assert RAM(8086) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8086)))) severity failure;
    assert RAM(8087) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8087)))) severity failure;
    assert RAM(8088) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8088)))) severity failure;
    assert RAM(8089) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8089)))) severity failure;
    assert RAM(8090) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8090)))) severity failure;
    assert RAM(8091) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8091)))) severity failure;
    assert RAM(8092) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8092)))) severity failure;
    assert RAM(8093) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8093)))) severity failure;
    assert RAM(8094) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8094)))) severity failure;
    assert RAM(8095) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8095)))) severity failure;
    assert RAM(8096) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8096)))) severity failure;
    assert RAM(8097) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8097)))) severity failure;
    assert RAM(8098) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8098)))) severity failure;
    assert RAM(8099) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8099)))) severity failure;
    assert RAM(8100) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8100)))) severity failure;
    assert RAM(8101) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8101)))) severity failure;
    assert RAM(8102) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8102)))) severity failure;
    assert RAM(8103) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8103)))) severity failure;
    assert RAM(8104) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8104)))) severity failure;
    assert RAM(8105) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8105)))) severity failure;
    assert RAM(8106) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8106)))) severity failure;
    assert RAM(8107) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8107)))) severity failure;
    assert RAM(8108) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8108)))) severity failure;
    assert RAM(8109) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8109)))) severity failure;
    assert RAM(8110) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8110)))) severity failure;
    assert RAM(8111) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8111)))) severity failure;
    assert RAM(8112) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8112)))) severity failure;
    assert RAM(8113) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8113)))) severity failure;
    assert RAM(8114) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8114)))) severity failure;
    assert RAM(8115) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8115)))) severity failure;
    assert RAM(8116) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8116)))) severity failure;
    assert RAM(8117) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8117)))) severity failure;
    assert RAM(8118) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8118)))) severity failure;
    assert RAM(8119) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8119)))) severity failure;
    assert RAM(8120) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8120)))) severity failure;
    assert RAM(8121) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8121)))) severity failure;
    assert RAM(8122) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8122)))) severity failure;
    assert RAM(8123) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8123)))) severity failure;
    assert RAM(8124) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8124)))) severity failure;
    assert RAM(8125) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8125)))) severity failure;
    assert RAM(8126) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8126)))) severity failure;
    assert RAM(8127) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8127)))) severity failure;
    assert RAM(8128) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8128)))) severity failure;
    assert RAM(8129) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8129)))) severity failure;
    assert RAM(8130) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8130)))) severity failure;
    assert RAM(8131) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8131)))) severity failure;
    assert RAM(8132) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8132)))) severity failure;
    assert RAM(8133) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8133)))) severity failure;
    assert RAM(8134) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8134)))) severity failure;
    assert RAM(8135) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8135)))) severity failure;
    assert RAM(8136) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8136)))) severity failure;
    assert RAM(8137) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8137)))) severity failure;
    assert RAM(8138) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8138)))) severity failure;
    assert RAM(8139) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8139)))) severity failure;
    assert RAM(8140) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8140)))) severity failure;
    assert RAM(8141) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8141)))) severity failure;
    assert RAM(8142) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8142)))) severity failure;
    assert RAM(8143) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8143)))) severity failure;
    assert RAM(8144) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8144)))) severity failure;
    assert RAM(8145) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8145)))) severity failure;
    assert RAM(8146) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8146)))) severity failure;
    assert RAM(8147) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8147)))) severity failure;
    assert RAM(8148) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8148)))) severity failure;
    assert RAM(8149) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8149)))) severity failure;
    assert RAM(8150) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8150)))) severity failure;
    assert RAM(8151) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8151)))) severity failure;
    assert RAM(8152) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8152)))) severity failure;
    assert RAM(8153) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8153)))) severity failure;
    assert RAM(8154) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8154)))) severity failure;
    assert RAM(8155) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8155)))) severity failure;
    assert RAM(8156) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8156)))) severity failure;
    assert RAM(8157) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8157)))) severity failure;
    assert RAM(8158) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8158)))) severity failure;
    assert RAM(8159) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8159)))) severity failure;
    assert RAM(8160) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8160)))) severity failure;
    assert RAM(8161) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8161)))) severity failure;
    assert RAM(8162) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8162)))) severity failure;
    assert RAM(8163) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8163)))) severity failure;
    assert RAM(8164) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8164)))) severity failure;
    assert RAM(8165) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8165)))) severity failure;
    assert RAM(8166) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8166)))) severity failure;
    assert RAM(8167) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8167)))) severity failure;
    assert RAM(8168) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8168)))) severity failure;
    assert RAM(8169) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8169)))) severity failure;
    assert RAM(8170) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8170)))) severity failure;
    assert RAM(8171) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8171)))) severity failure;
    assert RAM(8172) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8172)))) severity failure;
    assert RAM(8173) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8173)))) severity failure;
    assert RAM(8174) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8174)))) severity failure;
    assert RAM(8175) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8175)))) severity failure;
    assert RAM(8176) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8176)))) severity failure;
    assert RAM(8177) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8177)))) severity failure;
    assert RAM(8178) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8178)))) severity failure;
    assert RAM(8179) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8179)))) severity failure;
    assert RAM(8180) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8180)))) severity failure;
    assert RAM(8181) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8181)))) severity failure;
    assert RAM(8182) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8182)))) severity failure;
    assert RAM(8183) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8183)))) severity failure;
    assert RAM(8184) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8184)))) severity failure;
    assert RAM(8185) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8185)))) severity failure;
    assert RAM(8186) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8186)))) severity failure;
    assert RAM(8187) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8187)))) severity failure;
    assert RAM(8188) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8188)))) severity failure;
    assert RAM(8189) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8189)))) severity failure;
    assert RAM(8190) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8190)))) severity failure;
    assert RAM(8191) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8191)))) severity failure;
    assert RAM(8192) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8192)))) severity failure;
    assert RAM(8193) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8193)))) severity failure;
    assert RAM(8194) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8194)))) severity failure;
    assert RAM(8195) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8195)))) severity failure;
    assert RAM(8196) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8196)))) severity failure;
    assert RAM(8197) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8197)))) severity failure;
    assert RAM(8198) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8198)))) severity failure;
    assert RAM(8199) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8199)))) severity failure;
    assert RAM(8200) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8200)))) severity failure;
    assert RAM(8201) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8201)))) severity failure;
    assert RAM(8202) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8202)))) severity failure;
    assert RAM(8203) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8203)))) severity failure;
    assert RAM(8204) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8204)))) severity failure;
    assert RAM(8205) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8205)))) severity failure;
    assert RAM(8206) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8206)))) severity failure;
    assert RAM(8207) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8207)))) severity failure;
    assert RAM(8208) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8208)))) severity failure;
    assert RAM(8209) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8209)))) severity failure;
    assert RAM(8210) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8210)))) severity failure;
    assert RAM(8211) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8211)))) severity failure;
    assert RAM(8212) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8212)))) severity failure;
    assert RAM(8213) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8213)))) severity failure;
    assert RAM(8214) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8214)))) severity failure;
    assert RAM(8215) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8215)))) severity failure;
    assert RAM(8216) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8216)))) severity failure;
    assert RAM(8217) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8217)))) severity failure;
    assert RAM(8218) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8218)))) severity failure;
    assert RAM(8219) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8219)))) severity failure;
    assert RAM(8220) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8220)))) severity failure;
    assert RAM(8221) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8221)))) severity failure;
    assert RAM(8222) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8222)))) severity failure;
    assert RAM(8223) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8223)))) severity failure;
    assert RAM(8224) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8224)))) severity failure;
    assert RAM(8225) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8225)))) severity failure;
    assert RAM(8226) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8226)))) severity failure;
    assert RAM(8227) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8227)))) severity failure;
    assert RAM(8228) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8228)))) severity failure;
    assert RAM(8229) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8229)))) severity failure;
    assert RAM(8230) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8230)))) severity failure;
    assert RAM(8231) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8231)))) severity failure;
    assert RAM(8232) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8232)))) severity failure;
    assert RAM(8233) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8233)))) severity failure;
    assert RAM(8234) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8234)))) severity failure;
    assert RAM(8235) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8235)))) severity failure;
    assert RAM(8236) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8236)))) severity failure;
    assert RAM(8237) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8237)))) severity failure;
    assert RAM(8238) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8238)))) severity failure;
    assert RAM(8239) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8239)))) severity failure;
    assert RAM(8240) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8240)))) severity failure;
    assert RAM(8241) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8241)))) severity failure;
    assert RAM(8242) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8242)))) severity failure;
    assert RAM(8243) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8243)))) severity failure;
    assert RAM(8244) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8244)))) severity failure;
    assert RAM(8245) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8245)))) severity failure;
    assert RAM(8246) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8246)))) severity failure;
    assert RAM(8247) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8247)))) severity failure;
    assert RAM(8248) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8248)))) severity failure;
    assert RAM(8249) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8249)))) severity failure;
    assert RAM(8250) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8250)))) severity failure;
    assert RAM(8251) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8251)))) severity failure;
    assert RAM(8252) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8252)))) severity failure;
    assert RAM(8253) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8253)))) severity failure;
    assert RAM(8254) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8254)))) severity failure;
    assert RAM(8255) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8255)))) severity failure;
    assert RAM(8256) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8256)))) severity failure;
    assert RAM(8257) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8257)))) severity failure;
    assert RAM(8258) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8258)))) severity failure;
    assert RAM(8259) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8259)))) severity failure;
    assert RAM(8260) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8260)))) severity failure;
    assert RAM(8261) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8261)))) severity failure;
    assert RAM(8262) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8262)))) severity failure;
    assert RAM(8263) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8263)))) severity failure;
    assert RAM(8264) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8264)))) severity failure;
    assert RAM(8265) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8265)))) severity failure;
    assert RAM(8266) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8266)))) severity failure;
    assert RAM(8267) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8267)))) severity failure;
    assert RAM(8268) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8268)))) severity failure;
    assert RAM(8269) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8269)))) severity failure;
    assert RAM(8270) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8270)))) severity failure;
    assert RAM(8271) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8271)))) severity failure;
    assert RAM(8272) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8272)))) severity failure;
    assert RAM(8273) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8273)))) severity failure;
    assert RAM(8274) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8274)))) severity failure;
    assert RAM(8275) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8275)))) severity failure;
    assert RAM(8276) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8276)))) severity failure;
    assert RAM(8277) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8277)))) severity failure;
    assert RAM(8278) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8278)))) severity failure;
    assert RAM(8279) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8279)))) severity failure;
    assert RAM(8280) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8280)))) severity failure;
    assert RAM(8281) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8281)))) severity failure;
    assert RAM(8282) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8282)))) severity failure;
    assert RAM(8283) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8283)))) severity failure;
    assert RAM(8284) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8284)))) severity failure;
    assert RAM(8285) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8285)))) severity failure;
    assert RAM(8286) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8286)))) severity failure;
    assert RAM(8287) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8287)))) severity failure;
    assert RAM(8288) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8288)))) severity failure;
    assert RAM(8289) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8289)))) severity failure;
    assert RAM(8290) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8290)))) severity failure;
    assert RAM(8291) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8291)))) severity failure;
    assert RAM(8292) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8292)))) severity failure;
    assert RAM(8293) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8293)))) severity failure;
    assert RAM(8294) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8294)))) severity failure;
    assert RAM(8295) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8295)))) severity failure;
    assert RAM(8296) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8296)))) severity failure;
    assert RAM(8297) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8297)))) severity failure;
    assert RAM(8298) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8298)))) severity failure;
    assert RAM(8299) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8299)))) severity failure;
    assert RAM(8300) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8300)))) severity failure;
    assert RAM(8301) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8301)))) severity failure;
    assert RAM(8302) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8302)))) severity failure;
    assert RAM(8303) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8303)))) severity failure;
    assert RAM(8304) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8304)))) severity failure;
    assert RAM(8305) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8305)))) severity failure;
    assert RAM(8306) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8306)))) severity failure;
    assert RAM(8307) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8307)))) severity failure;
    assert RAM(8308) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8308)))) severity failure;
    assert RAM(8309) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8309)))) severity failure;
    assert RAM(8310) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8310)))) severity failure;
    assert RAM(8311) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8311)))) severity failure;
    assert RAM(8312) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8312)))) severity failure;
    assert RAM(8313) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8313)))) severity failure;
    assert RAM(8314) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8314)))) severity failure;
    assert RAM(8315) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8315)))) severity failure;
    assert RAM(8316) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8316)))) severity failure;
    assert RAM(8317) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8317)))) severity failure;
    assert RAM(8318) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8318)))) severity failure;
    assert RAM(8319) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8319)))) severity failure;
    assert RAM(8320) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8320)))) severity failure;
    assert RAM(8321) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8321)))) severity failure;
    assert RAM(8322) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8322)))) severity failure;
    assert RAM(8323) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8323)))) severity failure;
    assert RAM(8324) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8324)))) severity failure;
    assert RAM(8325) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8325)))) severity failure;
    assert RAM(8326) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8326)))) severity failure;
    assert RAM(8327) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8327)))) severity failure;
    assert RAM(8328) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8328)))) severity failure;
    assert RAM(8329) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8329)))) severity failure;
    assert RAM(8330) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8330)))) severity failure;
    assert RAM(8331) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8331)))) severity failure;
    assert RAM(8332) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8332)))) severity failure;
    assert RAM(8333) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8333)))) severity failure;
    assert RAM(8334) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8334)))) severity failure;
    assert RAM(8335) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8335)))) severity failure;
    assert RAM(8336) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8336)))) severity failure;
    assert RAM(8337) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8337)))) severity failure;
    assert RAM(8338) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8338)))) severity failure;
    assert RAM(8339) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8339)))) severity failure;
    assert RAM(8340) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8340)))) severity failure;
    assert RAM(8341) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8341)))) severity failure;
    assert RAM(8342) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8342)))) severity failure;
    assert RAM(8343) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8343)))) severity failure;
    assert RAM(8344) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8344)))) severity failure;
    assert RAM(8345) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8345)))) severity failure;
    assert RAM(8346) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8346)))) severity failure;
    assert RAM(8347) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(8347)))) severity failure;
    assert RAM(8348) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8348)))) severity failure;
    assert RAM(8349) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8349)))) severity failure;
    assert RAM(8350) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8350)))) severity failure;
    assert RAM(8351) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8351)))) severity failure;
    assert RAM(8352) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8352)))) severity failure;
    assert RAM(8353) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8353)))) severity failure;
    assert RAM(8354) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8354)))) severity failure;
    assert RAM(8355) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8355)))) severity failure;
    assert RAM(8356) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8356)))) severity failure;
    assert RAM(8357) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8357)))) severity failure;
    assert RAM(8358) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8358)))) severity failure;
    assert RAM(8359) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8359)))) severity failure;
    assert RAM(8360) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8360)))) severity failure;
    assert RAM(8361) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(8361)))) severity failure;
    assert RAM(8362) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(8362)))) severity failure;
    assert RAM(8363) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8363)))) severity failure;
    assert RAM(8364) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8364)))) severity failure;
    assert RAM(8365) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8365)))) severity failure;
    assert RAM(8366) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8366)))) severity failure;
    assert RAM(8367) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8367)))) severity failure;
    assert RAM(8368) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8368)))) severity failure;
    assert RAM(8369) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8369)))) severity failure;
    assert RAM(8370) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8370)))) severity failure;
    assert RAM(8371) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8371)))) severity failure;
    assert RAM(8372) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8372)))) severity failure;
    assert RAM(8373) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8373)))) severity failure;
    assert RAM(8374) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(8374)))) severity failure;
    assert RAM(8375) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(8375)))) severity failure;
    assert RAM(8376) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8376)))) severity failure;
    assert RAM(8377) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8377)))) severity failure;
    assert RAM(8378) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(8378)))) severity failure;
    assert RAM(8379) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(8379)))) severity failure;

    assert false report "Simulation Ended! TEST PASSATO" severity failure;
end process test;

end shlev5tb;
