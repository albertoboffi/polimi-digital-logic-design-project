-------------------------------------------------------------------------------
--
-- Final examination - Digital Logic Design
-- Alberto Boffi - Politecnico di Milano, AY 2020/21
-- TEST MODULE: Shift level = 7
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity shlev7_tb is
end shlev7_tb;

architecture shlev7tb of shlev7_tb is
constant c_CLOCK_PERIOD         : time := 15 ns;
signal   tb_done                : std_logic;
signal   mem_address            : std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst                 : std_logic := '0';
signal   tb_start               : std_logic := '0';
signal   tb_clk                 : std_logic := '0';
signal   mem_o_data,mem_i_data  : std_logic_vector (7 downto 0);
signal   enable_wire            : std_logic;
signal   mem_we                 : std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);


signal RAM: ram_type :=
	(0 => std_logic_vector(to_unsigned(73, 8)),
	1 => std_logic_vector(to_unsigned(92, 8)),
	2 => std_logic_vector(to_unsigned(41, 8)),
	3 => std_logic_vector(to_unsigned(41, 8)),
	4 => std_logic_vector(to_unsigned(42, 8)),
	5 => std_logic_vector(to_unsigned(42, 8)),
	6 => std_logic_vector(to_unsigned(42, 8)),
	7 => std_logic_vector(to_unsigned(41, 8)),
	8 => std_logic_vector(to_unsigned(41, 8)),
	9 => std_logic_vector(to_unsigned(41, 8)),
	10 => std_logic_vector(to_unsigned(41, 8)),
	11 => std_logic_vector(to_unsigned(42, 8)),
	12 => std_logic_vector(to_unsigned(41, 8)),
	13 => std_logic_vector(to_unsigned(42, 8)),
	14 => std_logic_vector(to_unsigned(42, 8)),
	15 => std_logic_vector(to_unsigned(41, 8)),
	16 => std_logic_vector(to_unsigned(42, 8)),
	17 => std_logic_vector(to_unsigned(42, 8)),
	18 => std_logic_vector(to_unsigned(42, 8)),
	19 => std_logic_vector(to_unsigned(41, 8)),
	20 => std_logic_vector(to_unsigned(42, 8)),
	21 => std_logic_vector(to_unsigned(41, 8)),
	22 => std_logic_vector(to_unsigned(41, 8)),
	23 => std_logic_vector(to_unsigned(41, 8)),
	24 => std_logic_vector(to_unsigned(42, 8)),
	25 => std_logic_vector(to_unsigned(41, 8)),
	26 => std_logic_vector(to_unsigned(42, 8)),
	27 => std_logic_vector(to_unsigned(41, 8)),
	28 => std_logic_vector(to_unsigned(41, 8)),
	29 => std_logic_vector(to_unsigned(41, 8)),
	30 => std_logic_vector(to_unsigned(42, 8)),
	31 => std_logic_vector(to_unsigned(42, 8)),
	32 => std_logic_vector(to_unsigned(42, 8)),
	33 => std_logic_vector(to_unsigned(42, 8)),
	34 => std_logic_vector(to_unsigned(42, 8)),
	35 => std_logic_vector(to_unsigned(42, 8)),
	36 => std_logic_vector(to_unsigned(41, 8)),
	37 => std_logic_vector(to_unsigned(41, 8)),
	38 => std_logic_vector(to_unsigned(41, 8)),
	39 => std_logic_vector(to_unsigned(42, 8)),
	40 => std_logic_vector(to_unsigned(41, 8)),
	41 => std_logic_vector(to_unsigned(41, 8)),
	42 => std_logic_vector(to_unsigned(42, 8)),
	43 => std_logic_vector(to_unsigned(42, 8)),
	44 => std_logic_vector(to_unsigned(42, 8)),
	45 => std_logic_vector(to_unsigned(41, 8)),
	46 => std_logic_vector(to_unsigned(41, 8)),
	47 => std_logic_vector(to_unsigned(42, 8)),
	48 => std_logic_vector(to_unsigned(42, 8)),
	49 => std_logic_vector(to_unsigned(42, 8)),
	50 => std_logic_vector(to_unsigned(41, 8)),
	51 => std_logic_vector(to_unsigned(42, 8)),
	52 => std_logic_vector(to_unsigned(42, 8)),
	53 => std_logic_vector(to_unsigned(42, 8)),
	54 => std_logic_vector(to_unsigned(41, 8)),
	55 => std_logic_vector(to_unsigned(41, 8)),
	56 => std_logic_vector(to_unsigned(41, 8)),
	57 => std_logic_vector(to_unsigned(41, 8)),
	58 => std_logic_vector(to_unsigned(41, 8)),
	59 => std_logic_vector(to_unsigned(41, 8)),
	60 => std_logic_vector(to_unsigned(42, 8)),
	61 => std_logic_vector(to_unsigned(42, 8)),
	62 => std_logic_vector(to_unsigned(41, 8)),
	63 => std_logic_vector(to_unsigned(41, 8)),
	64 => std_logic_vector(to_unsigned(42, 8)),
	65 => std_logic_vector(to_unsigned(41, 8)),
	66 => std_logic_vector(to_unsigned(42, 8)),
	67 => std_logic_vector(to_unsigned(42, 8)),
	68 => std_logic_vector(to_unsigned(41, 8)),
	69 => std_logic_vector(to_unsigned(41, 8)),
	70 => std_logic_vector(to_unsigned(42, 8)),
	71 => std_logic_vector(to_unsigned(42, 8)),
	72 => std_logic_vector(to_unsigned(42, 8)),
	73 => std_logic_vector(to_unsigned(41, 8)),
	74 => std_logic_vector(to_unsigned(42, 8)),
	75 => std_logic_vector(to_unsigned(42, 8)),
	76 => std_logic_vector(to_unsigned(41, 8)),
	77 => std_logic_vector(to_unsigned(41, 8)),
	78 => std_logic_vector(to_unsigned(42, 8)),
	79 => std_logic_vector(to_unsigned(42, 8)),
	80 => std_logic_vector(to_unsigned(42, 8)),
	81 => std_logic_vector(to_unsigned(41, 8)),
	82 => std_logic_vector(to_unsigned(41, 8)),
	83 => std_logic_vector(to_unsigned(42, 8)),
	84 => std_logic_vector(to_unsigned(41, 8)),
	85 => std_logic_vector(to_unsigned(42, 8)),
	86 => std_logic_vector(to_unsigned(41, 8)),
	87 => std_logic_vector(to_unsigned(41, 8)),
	88 => std_logic_vector(to_unsigned(42, 8)),
	89 => std_logic_vector(to_unsigned(42, 8)),
	90 => std_logic_vector(to_unsigned(42, 8)),
	91 => std_logic_vector(to_unsigned(42, 8)),
	92 => std_logic_vector(to_unsigned(41, 8)),
	93 => std_logic_vector(to_unsigned(42, 8)),
	94 => std_logic_vector(to_unsigned(42, 8)),
	95 => std_logic_vector(to_unsigned(41, 8)),
	96 => std_logic_vector(to_unsigned(41, 8)),
	97 => std_logic_vector(to_unsigned(42, 8)),
	98 => std_logic_vector(to_unsigned(41, 8)),
	99 => std_logic_vector(to_unsigned(41, 8)),
	100 => std_logic_vector(to_unsigned(42, 8)),
	101 => std_logic_vector(to_unsigned(41, 8)),
	102 => std_logic_vector(to_unsigned(42, 8)),
	103 => std_logic_vector(to_unsigned(42, 8)),
	104 => std_logic_vector(to_unsigned(41, 8)),
	105 => std_logic_vector(to_unsigned(42, 8)),
	106 => std_logic_vector(to_unsigned(42, 8)),
	107 => std_logic_vector(to_unsigned(42, 8)),
	108 => std_logic_vector(to_unsigned(42, 8)),
	109 => std_logic_vector(to_unsigned(41, 8)),
	110 => std_logic_vector(to_unsigned(41, 8)),
	111 => std_logic_vector(to_unsigned(41, 8)),
	112 => std_logic_vector(to_unsigned(42, 8)),
	113 => std_logic_vector(to_unsigned(41, 8)),
	114 => std_logic_vector(to_unsigned(42, 8)),
	115 => std_logic_vector(to_unsigned(41, 8)),
	116 => std_logic_vector(to_unsigned(42, 8)),
	117 => std_logic_vector(to_unsigned(42, 8)),
	118 => std_logic_vector(to_unsigned(41, 8)),
	119 => std_logic_vector(to_unsigned(41, 8)),
	120 => std_logic_vector(to_unsigned(41, 8)),
	121 => std_logic_vector(to_unsigned(42, 8)),
	122 => std_logic_vector(to_unsigned(41, 8)),
	123 => std_logic_vector(to_unsigned(41, 8)),
	124 => std_logic_vector(to_unsigned(42, 8)),
	125 => std_logic_vector(to_unsigned(42, 8)),
	126 => std_logic_vector(to_unsigned(41, 8)),
	127 => std_logic_vector(to_unsigned(41, 8)),
	128 => std_logic_vector(to_unsigned(41, 8)),
	129 => std_logic_vector(to_unsigned(42, 8)),
	130 => std_logic_vector(to_unsigned(42, 8)),
	131 => std_logic_vector(to_unsigned(42, 8)),
	132 => std_logic_vector(to_unsigned(42, 8)),
	133 => std_logic_vector(to_unsigned(42, 8)),
	134 => std_logic_vector(to_unsigned(41, 8)),
	135 => std_logic_vector(to_unsigned(42, 8)),
	136 => std_logic_vector(to_unsigned(41, 8)),
	137 => std_logic_vector(to_unsigned(42, 8)),
	138 => std_logic_vector(to_unsigned(41, 8)),
	139 => std_logic_vector(to_unsigned(41, 8)),
	140 => std_logic_vector(to_unsigned(41, 8)),
	141 => std_logic_vector(to_unsigned(41, 8)),
	142 => std_logic_vector(to_unsigned(42, 8)),
	143 => std_logic_vector(to_unsigned(42, 8)),
	144 => std_logic_vector(to_unsigned(42, 8)),
	145 => std_logic_vector(to_unsigned(42, 8)),
	146 => std_logic_vector(to_unsigned(42, 8)),
	147 => std_logic_vector(to_unsigned(41, 8)),
	148 => std_logic_vector(to_unsigned(42, 8)),
	149 => std_logic_vector(to_unsigned(42, 8)),
	150 => std_logic_vector(to_unsigned(41, 8)),
	151 => std_logic_vector(to_unsigned(41, 8)),
	152 => std_logic_vector(to_unsigned(41, 8)),
	153 => std_logic_vector(to_unsigned(42, 8)),
	154 => std_logic_vector(to_unsigned(42, 8)),
	155 => std_logic_vector(to_unsigned(41, 8)),
	156 => std_logic_vector(to_unsigned(42, 8)),
	157 => std_logic_vector(to_unsigned(42, 8)),
	158 => std_logic_vector(to_unsigned(41, 8)),
	159 => std_logic_vector(to_unsigned(41, 8)),
	160 => std_logic_vector(to_unsigned(41, 8)),
	161 => std_logic_vector(to_unsigned(42, 8)),
	162 => std_logic_vector(to_unsigned(41, 8)),
	163 => std_logic_vector(to_unsigned(41, 8)),
	164 => std_logic_vector(to_unsigned(41, 8)),
	165 => std_logic_vector(to_unsigned(42, 8)),
	166 => std_logic_vector(to_unsigned(42, 8)),
	167 => std_logic_vector(to_unsigned(42, 8)),
	168 => std_logic_vector(to_unsigned(41, 8)),
	169 => std_logic_vector(to_unsigned(42, 8)),
	170 => std_logic_vector(to_unsigned(42, 8)),
	171 => std_logic_vector(to_unsigned(41, 8)),
	172 => std_logic_vector(to_unsigned(42, 8)),
	173 => std_logic_vector(to_unsigned(42, 8)),
	174 => std_logic_vector(to_unsigned(41, 8)),
	175 => std_logic_vector(to_unsigned(41, 8)),
	176 => std_logic_vector(to_unsigned(42, 8)),
	177 => std_logic_vector(to_unsigned(42, 8)),
	178 => std_logic_vector(to_unsigned(42, 8)),
	179 => std_logic_vector(to_unsigned(41, 8)),
	180 => std_logic_vector(to_unsigned(42, 8)),
	181 => std_logic_vector(to_unsigned(41, 8)),
	182 => std_logic_vector(to_unsigned(42, 8)),
	183 => std_logic_vector(to_unsigned(41, 8)),
	184 => std_logic_vector(to_unsigned(42, 8)),
	185 => std_logic_vector(to_unsigned(41, 8)),
	186 => std_logic_vector(to_unsigned(42, 8)),
	187 => std_logic_vector(to_unsigned(42, 8)),
	188 => std_logic_vector(to_unsigned(41, 8)),
	189 => std_logic_vector(to_unsigned(41, 8)),
	190 => std_logic_vector(to_unsigned(42, 8)),
	191 => std_logic_vector(to_unsigned(42, 8)),
	192 => std_logic_vector(to_unsigned(42, 8)),
	193 => std_logic_vector(to_unsigned(42, 8)),
	194 => std_logic_vector(to_unsigned(41, 8)),
	195 => std_logic_vector(to_unsigned(41, 8)),
	196 => std_logic_vector(to_unsigned(42, 8)),
	197 => std_logic_vector(to_unsigned(41, 8)),
	198 => std_logic_vector(to_unsigned(42, 8)),
	199 => std_logic_vector(to_unsigned(41, 8)),
	200 => std_logic_vector(to_unsigned(42, 8)),
	201 => std_logic_vector(to_unsigned(42, 8)),
	202 => std_logic_vector(to_unsigned(41, 8)),
	203 => std_logic_vector(to_unsigned(41, 8)),
	204 => std_logic_vector(to_unsigned(41, 8)),
	205 => std_logic_vector(to_unsigned(41, 8)),
	206 => std_logic_vector(to_unsigned(42, 8)),
	207 => std_logic_vector(to_unsigned(41, 8)),
	208 => std_logic_vector(to_unsigned(41, 8)),
	209 => std_logic_vector(to_unsigned(42, 8)),
	210 => std_logic_vector(to_unsigned(41, 8)),
	211 => std_logic_vector(to_unsigned(41, 8)),
	212 => std_logic_vector(to_unsigned(42, 8)),
	213 => std_logic_vector(to_unsigned(42, 8)),
	214 => std_logic_vector(to_unsigned(42, 8)),
	215 => std_logic_vector(to_unsigned(41, 8)),
	216 => std_logic_vector(to_unsigned(42, 8)),
	217 => std_logic_vector(to_unsigned(42, 8)),
	218 => std_logic_vector(to_unsigned(41, 8)),
	219 => std_logic_vector(to_unsigned(41, 8)),
	220 => std_logic_vector(to_unsigned(41, 8)),
	221 => std_logic_vector(to_unsigned(41, 8)),
	222 => std_logic_vector(to_unsigned(42, 8)),
	223 => std_logic_vector(to_unsigned(42, 8)),
	224 => std_logic_vector(to_unsigned(42, 8)),
	225 => std_logic_vector(to_unsigned(41, 8)),
	226 => std_logic_vector(to_unsigned(41, 8)),
	227 => std_logic_vector(to_unsigned(42, 8)),
	228 => std_logic_vector(to_unsigned(42, 8)),
	229 => std_logic_vector(to_unsigned(42, 8)),
	230 => std_logic_vector(to_unsigned(42, 8)),
	231 => std_logic_vector(to_unsigned(42, 8)),
	232 => std_logic_vector(to_unsigned(42, 8)),
	233 => std_logic_vector(to_unsigned(41, 8)),
	234 => std_logic_vector(to_unsigned(41, 8)),
	235 => std_logic_vector(to_unsigned(42, 8)),
	236 => std_logic_vector(to_unsigned(42, 8)),
	237 => std_logic_vector(to_unsigned(41, 8)),
	238 => std_logic_vector(to_unsigned(42, 8)),
	239 => std_logic_vector(to_unsigned(41, 8)),
	240 => std_logic_vector(to_unsigned(41, 8)),
	241 => std_logic_vector(to_unsigned(41, 8)),
	242 => std_logic_vector(to_unsigned(42, 8)),
	243 => std_logic_vector(to_unsigned(41, 8)),
	244 => std_logic_vector(to_unsigned(42, 8)),
	245 => std_logic_vector(to_unsigned(42, 8)),
	246 => std_logic_vector(to_unsigned(42, 8)),
	247 => std_logic_vector(to_unsigned(41, 8)),
	248 => std_logic_vector(to_unsigned(41, 8)),
	249 => std_logic_vector(to_unsigned(42, 8)),
	250 => std_logic_vector(to_unsigned(42, 8)),
	251 => std_logic_vector(to_unsigned(41, 8)),
	252 => std_logic_vector(to_unsigned(42, 8)),
	253 => std_logic_vector(to_unsigned(41, 8)),
	254 => std_logic_vector(to_unsigned(41, 8)),
	255 => std_logic_vector(to_unsigned(41, 8)),
	256 => std_logic_vector(to_unsigned(41, 8)),
	257 => std_logic_vector(to_unsigned(41, 8)),
	258 => std_logic_vector(to_unsigned(42, 8)),
	259 => std_logic_vector(to_unsigned(41, 8)),
	260 => std_logic_vector(to_unsigned(42, 8)),
	261 => std_logic_vector(to_unsigned(42, 8)),
	262 => std_logic_vector(to_unsigned(42, 8)),
	263 => std_logic_vector(to_unsigned(41, 8)),
	264 => std_logic_vector(to_unsigned(41, 8)),
	265 => std_logic_vector(to_unsigned(42, 8)),
	266 => std_logic_vector(to_unsigned(42, 8)),
	267 => std_logic_vector(to_unsigned(41, 8)),
	268 => std_logic_vector(to_unsigned(42, 8)),
	269 => std_logic_vector(to_unsigned(41, 8)),
	270 => std_logic_vector(to_unsigned(42, 8)),
	271 => std_logic_vector(to_unsigned(42, 8)),
	272 => std_logic_vector(to_unsigned(42, 8)),
	273 => std_logic_vector(to_unsigned(41, 8)),
	274 => std_logic_vector(to_unsigned(41, 8)),
	275 => std_logic_vector(to_unsigned(42, 8)),
	276 => std_logic_vector(to_unsigned(41, 8)),
	277 => std_logic_vector(to_unsigned(42, 8)),
	278 => std_logic_vector(to_unsigned(42, 8)),
	279 => std_logic_vector(to_unsigned(42, 8)),
	280 => std_logic_vector(to_unsigned(42, 8)),
	281 => std_logic_vector(to_unsigned(42, 8)),
	282 => std_logic_vector(to_unsigned(42, 8)),
	283 => std_logic_vector(to_unsigned(42, 8)),
	284 => std_logic_vector(to_unsigned(41, 8)),
	285 => std_logic_vector(to_unsigned(42, 8)),
	286 => std_logic_vector(to_unsigned(42, 8)),
	287 => std_logic_vector(to_unsigned(42, 8)),
	288 => std_logic_vector(to_unsigned(41, 8)),
	289 => std_logic_vector(to_unsigned(42, 8)),
	290 => std_logic_vector(to_unsigned(41, 8)),
	291 => std_logic_vector(to_unsigned(42, 8)),
	292 => std_logic_vector(to_unsigned(42, 8)),
	293 => std_logic_vector(to_unsigned(41, 8)),
	294 => std_logic_vector(to_unsigned(42, 8)),
	295 => std_logic_vector(to_unsigned(42, 8)),
	296 => std_logic_vector(to_unsigned(41, 8)),
	297 => std_logic_vector(to_unsigned(41, 8)),
	298 => std_logic_vector(to_unsigned(42, 8)),
	299 => std_logic_vector(to_unsigned(41, 8)),
	300 => std_logic_vector(to_unsigned(42, 8)),
	301 => std_logic_vector(to_unsigned(42, 8)),
	302 => std_logic_vector(to_unsigned(42, 8)),
	303 => std_logic_vector(to_unsigned(42, 8)),
	304 => std_logic_vector(to_unsigned(42, 8)),
	305 => std_logic_vector(to_unsigned(41, 8)),
	306 => std_logic_vector(to_unsigned(41, 8)),
	307 => std_logic_vector(to_unsigned(42, 8)),
	308 => std_logic_vector(to_unsigned(42, 8)),
	309 => std_logic_vector(to_unsigned(42, 8)),
	310 => std_logic_vector(to_unsigned(41, 8)),
	311 => std_logic_vector(to_unsigned(41, 8)),
	312 => std_logic_vector(to_unsigned(42, 8)),
	313 => std_logic_vector(to_unsigned(41, 8)),
	314 => std_logic_vector(to_unsigned(41, 8)),
	315 => std_logic_vector(to_unsigned(41, 8)),
	316 => std_logic_vector(to_unsigned(41, 8)),
	317 => std_logic_vector(to_unsigned(41, 8)),
	318 => std_logic_vector(to_unsigned(42, 8)),
	319 => std_logic_vector(to_unsigned(41, 8)),
	320 => std_logic_vector(to_unsigned(41, 8)),
	321 => std_logic_vector(to_unsigned(41, 8)),
	322 => std_logic_vector(to_unsigned(41, 8)),
	323 => std_logic_vector(to_unsigned(41, 8)),
	324 => std_logic_vector(to_unsigned(41, 8)),
	325 => std_logic_vector(to_unsigned(42, 8)),
	326 => std_logic_vector(to_unsigned(42, 8)),
	327 => std_logic_vector(to_unsigned(42, 8)),
	328 => std_logic_vector(to_unsigned(42, 8)),
	329 => std_logic_vector(to_unsigned(41, 8)),
	330 => std_logic_vector(to_unsigned(42, 8)),
	331 => std_logic_vector(to_unsigned(41, 8)),
	332 => std_logic_vector(to_unsigned(42, 8)),
	333 => std_logic_vector(to_unsigned(42, 8)),
	334 => std_logic_vector(to_unsigned(42, 8)),
	335 => std_logic_vector(to_unsigned(42, 8)),
	336 => std_logic_vector(to_unsigned(41, 8)),
	337 => std_logic_vector(to_unsigned(41, 8)),
	338 => std_logic_vector(to_unsigned(41, 8)),
	339 => std_logic_vector(to_unsigned(42, 8)),
	340 => std_logic_vector(to_unsigned(42, 8)),
	341 => std_logic_vector(to_unsigned(41, 8)),
	342 => std_logic_vector(to_unsigned(42, 8)),
	343 => std_logic_vector(to_unsigned(42, 8)),
	344 => std_logic_vector(to_unsigned(41, 8)),
	345 => std_logic_vector(to_unsigned(41, 8)),
	346 => std_logic_vector(to_unsigned(41, 8)),
	347 => std_logic_vector(to_unsigned(42, 8)),
	348 => std_logic_vector(to_unsigned(42, 8)),
	349 => std_logic_vector(to_unsigned(41, 8)),
	350 => std_logic_vector(to_unsigned(41, 8)),
	351 => std_logic_vector(to_unsigned(41, 8)),
	352 => std_logic_vector(to_unsigned(42, 8)),
	353 => std_logic_vector(to_unsigned(41, 8)),
	354 => std_logic_vector(to_unsigned(41, 8)),
	355 => std_logic_vector(to_unsigned(41, 8)),
	356 => std_logic_vector(to_unsigned(41, 8)),
	357 => std_logic_vector(to_unsigned(41, 8)),
	358 => std_logic_vector(to_unsigned(41, 8)),
	359 => std_logic_vector(to_unsigned(41, 8)),
	360 => std_logic_vector(to_unsigned(41, 8)),
	361 => std_logic_vector(to_unsigned(41, 8)),
	362 => std_logic_vector(to_unsigned(42, 8)),
	363 => std_logic_vector(to_unsigned(42, 8)),
	364 => std_logic_vector(to_unsigned(41, 8)),
	365 => std_logic_vector(to_unsigned(42, 8)),
	366 => std_logic_vector(to_unsigned(42, 8)),
	367 => std_logic_vector(to_unsigned(42, 8)),
	368 => std_logic_vector(to_unsigned(42, 8)),
	369 => std_logic_vector(to_unsigned(41, 8)),
	370 => std_logic_vector(to_unsigned(41, 8)),
	371 => std_logic_vector(to_unsigned(41, 8)),
	372 => std_logic_vector(to_unsigned(42, 8)),
	373 => std_logic_vector(to_unsigned(42, 8)),
	374 => std_logic_vector(to_unsigned(41, 8)),
	375 => std_logic_vector(to_unsigned(42, 8)),
	376 => std_logic_vector(to_unsigned(42, 8)),
	377 => std_logic_vector(to_unsigned(41, 8)),
	378 => std_logic_vector(to_unsigned(41, 8)),
	379 => std_logic_vector(to_unsigned(41, 8)),
	380 => std_logic_vector(to_unsigned(42, 8)),
	381 => std_logic_vector(to_unsigned(41, 8)),
	382 => std_logic_vector(to_unsigned(41, 8)),
	383 => std_logic_vector(to_unsigned(42, 8)),
	384 => std_logic_vector(to_unsigned(41, 8)),
	385 => std_logic_vector(to_unsigned(41, 8)),
	386 => std_logic_vector(to_unsigned(41, 8)),
	387 => std_logic_vector(to_unsigned(41, 8)),
	388 => std_logic_vector(to_unsigned(42, 8)),
	389 => std_logic_vector(to_unsigned(42, 8)),
	390 => std_logic_vector(to_unsigned(42, 8)),
	391 => std_logic_vector(to_unsigned(42, 8)),
	392 => std_logic_vector(to_unsigned(41, 8)),
	393 => std_logic_vector(to_unsigned(41, 8)),
	394 => std_logic_vector(to_unsigned(42, 8)),
	395 => std_logic_vector(to_unsigned(42, 8)),
	396 => std_logic_vector(to_unsigned(42, 8)),
	397 => std_logic_vector(to_unsigned(41, 8)),
	398 => std_logic_vector(to_unsigned(41, 8)),
	399 => std_logic_vector(to_unsigned(42, 8)),
	400 => std_logic_vector(to_unsigned(41, 8)),
	401 => std_logic_vector(to_unsigned(41, 8)),
	402 => std_logic_vector(to_unsigned(41, 8)),
	403 => std_logic_vector(to_unsigned(41, 8)),
	404 => std_logic_vector(to_unsigned(41, 8)),
	405 => std_logic_vector(to_unsigned(42, 8)),
	406 => std_logic_vector(to_unsigned(41, 8)),
	407 => std_logic_vector(to_unsigned(41, 8)),
	408 => std_logic_vector(to_unsigned(42, 8)),
	409 => std_logic_vector(to_unsigned(42, 8)),
	410 => std_logic_vector(to_unsigned(42, 8)),
	411 => std_logic_vector(to_unsigned(41, 8)),
	412 => std_logic_vector(to_unsigned(42, 8)),
	413 => std_logic_vector(to_unsigned(42, 8)),
	414 => std_logic_vector(to_unsigned(42, 8)),
	415 => std_logic_vector(to_unsigned(42, 8)),
	416 => std_logic_vector(to_unsigned(41, 8)),
	417 => std_logic_vector(to_unsigned(41, 8)),
	418 => std_logic_vector(to_unsigned(41, 8)),
	419 => std_logic_vector(to_unsigned(41, 8)),
	420 => std_logic_vector(to_unsigned(42, 8)),
	421 => std_logic_vector(to_unsigned(41, 8)),
	422 => std_logic_vector(to_unsigned(42, 8)),
	423 => std_logic_vector(to_unsigned(41, 8)),
	424 => std_logic_vector(to_unsigned(41, 8)),
	425 => std_logic_vector(to_unsigned(41, 8)),
	426 => std_logic_vector(to_unsigned(42, 8)),
	427 => std_logic_vector(to_unsigned(42, 8)),
	428 => std_logic_vector(to_unsigned(42, 8)),
	429 => std_logic_vector(to_unsigned(42, 8)),
	430 => std_logic_vector(to_unsigned(42, 8)),
	431 => std_logic_vector(to_unsigned(42, 8)),
	432 => std_logic_vector(to_unsigned(41, 8)),
	433 => std_logic_vector(to_unsigned(42, 8)),
	434 => std_logic_vector(to_unsigned(41, 8)),
	435 => std_logic_vector(to_unsigned(42, 8)),
	436 => std_logic_vector(to_unsigned(41, 8)),
	437 => std_logic_vector(to_unsigned(41, 8)),
	438 => std_logic_vector(to_unsigned(41, 8)),
	439 => std_logic_vector(to_unsigned(41, 8)),
	440 => std_logic_vector(to_unsigned(41, 8)),
	441 => std_logic_vector(to_unsigned(41, 8)),
	442 => std_logic_vector(to_unsigned(42, 8)),
	443 => std_logic_vector(to_unsigned(42, 8)),
	444 => std_logic_vector(to_unsigned(42, 8)),
	445 => std_logic_vector(to_unsigned(42, 8)),
	446 => std_logic_vector(to_unsigned(41, 8)),
	447 => std_logic_vector(to_unsigned(42, 8)),
	448 => std_logic_vector(to_unsigned(42, 8)),
	449 => std_logic_vector(to_unsigned(41, 8)),
	450 => std_logic_vector(to_unsigned(42, 8)),
	451 => std_logic_vector(to_unsigned(41, 8)),
	452 => std_logic_vector(to_unsigned(42, 8)),
	453 => std_logic_vector(to_unsigned(42, 8)),
	454 => std_logic_vector(to_unsigned(42, 8)),
	455 => std_logic_vector(to_unsigned(42, 8)),
	456 => std_logic_vector(to_unsigned(41, 8)),
	457 => std_logic_vector(to_unsigned(41, 8)),
	458 => std_logic_vector(to_unsigned(41, 8)),
	459 => std_logic_vector(to_unsigned(42, 8)),
	460 => std_logic_vector(to_unsigned(42, 8)),
	461 => std_logic_vector(to_unsigned(41, 8)),
	462 => std_logic_vector(to_unsigned(41, 8)),
	463 => std_logic_vector(to_unsigned(41, 8)),
	464 => std_logic_vector(to_unsigned(41, 8)),
	465 => std_logic_vector(to_unsigned(41, 8)),
	466 => std_logic_vector(to_unsigned(41, 8)),
	467 => std_logic_vector(to_unsigned(42, 8)),
	468 => std_logic_vector(to_unsigned(41, 8)),
	469 => std_logic_vector(to_unsigned(41, 8)),
	470 => std_logic_vector(to_unsigned(41, 8)),
	471 => std_logic_vector(to_unsigned(41, 8)),
	472 => std_logic_vector(to_unsigned(41, 8)),
	473 => std_logic_vector(to_unsigned(41, 8)),
	474 => std_logic_vector(to_unsigned(42, 8)),
	475 => std_logic_vector(to_unsigned(41, 8)),
	476 => std_logic_vector(to_unsigned(41, 8)),
	477 => std_logic_vector(to_unsigned(41, 8)),
	478 => std_logic_vector(to_unsigned(41, 8)),
	479 => std_logic_vector(to_unsigned(42, 8)),
	480 => std_logic_vector(to_unsigned(41, 8)),
	481 => std_logic_vector(to_unsigned(41, 8)),
	482 => std_logic_vector(to_unsigned(42, 8)),
	483 => std_logic_vector(to_unsigned(42, 8)),
	484 => std_logic_vector(to_unsigned(42, 8)),
	485 => std_logic_vector(to_unsigned(41, 8)),
	486 => std_logic_vector(to_unsigned(41, 8)),
	487 => std_logic_vector(to_unsigned(41, 8)),
	488 => std_logic_vector(to_unsigned(41, 8)),
	489 => std_logic_vector(to_unsigned(41, 8)),
	490 => std_logic_vector(to_unsigned(42, 8)),
	491 => std_logic_vector(to_unsigned(42, 8)),
	492 => std_logic_vector(to_unsigned(41, 8)),
	493 => std_logic_vector(to_unsigned(41, 8)),
	494 => std_logic_vector(to_unsigned(42, 8)),
	495 => std_logic_vector(to_unsigned(41, 8)),
	496 => std_logic_vector(to_unsigned(41, 8)),
	497 => std_logic_vector(to_unsigned(42, 8)),
	498 => std_logic_vector(to_unsigned(41, 8)),
	499 => std_logic_vector(to_unsigned(41, 8)),
	500 => std_logic_vector(to_unsigned(42, 8)),
	501 => std_logic_vector(to_unsigned(41, 8)),
	502 => std_logic_vector(to_unsigned(41, 8)),
	503 => std_logic_vector(to_unsigned(42, 8)),
	504 => std_logic_vector(to_unsigned(42, 8)),
	505 => std_logic_vector(to_unsigned(41, 8)),
	506 => std_logic_vector(to_unsigned(41, 8)),
	507 => std_logic_vector(to_unsigned(42, 8)),
	508 => std_logic_vector(to_unsigned(42, 8)),
	509 => std_logic_vector(to_unsigned(42, 8)),
	510 => std_logic_vector(to_unsigned(42, 8)),
	511 => std_logic_vector(to_unsigned(42, 8)),
	512 => std_logic_vector(to_unsigned(41, 8)),
	513 => std_logic_vector(to_unsigned(41, 8)),
	514 => std_logic_vector(to_unsigned(42, 8)),
	515 => std_logic_vector(to_unsigned(42, 8)),
	516 => std_logic_vector(to_unsigned(41, 8)),
	517 => std_logic_vector(to_unsigned(42, 8)),
	518 => std_logic_vector(to_unsigned(41, 8)),
	519 => std_logic_vector(to_unsigned(42, 8)),
	520 => std_logic_vector(to_unsigned(41, 8)),
	521 => std_logic_vector(to_unsigned(42, 8)),
	522 => std_logic_vector(to_unsigned(41, 8)),
	523 => std_logic_vector(to_unsigned(42, 8)),
	524 => std_logic_vector(to_unsigned(42, 8)),
	525 => std_logic_vector(to_unsigned(41, 8)),
	526 => std_logic_vector(to_unsigned(42, 8)),
	527 => std_logic_vector(to_unsigned(41, 8)),
	528 => std_logic_vector(to_unsigned(42, 8)),
	529 => std_logic_vector(to_unsigned(42, 8)),
	530 => std_logic_vector(to_unsigned(42, 8)),
	531 => std_logic_vector(to_unsigned(42, 8)),
	532 => std_logic_vector(to_unsigned(41, 8)),
	533 => std_logic_vector(to_unsigned(42, 8)),
	534 => std_logic_vector(to_unsigned(42, 8)),
	535 => std_logic_vector(to_unsigned(42, 8)),
	536 => std_logic_vector(to_unsigned(41, 8)),
	537 => std_logic_vector(to_unsigned(42, 8)),
	538 => std_logic_vector(to_unsigned(42, 8)),
	539 => std_logic_vector(to_unsigned(41, 8)),
	540 => std_logic_vector(to_unsigned(42, 8)),
	541 => std_logic_vector(to_unsigned(42, 8)),
	542 => std_logic_vector(to_unsigned(42, 8)),
	543 => std_logic_vector(to_unsigned(41, 8)),
	544 => std_logic_vector(to_unsigned(41, 8)),
	545 => std_logic_vector(to_unsigned(41, 8)),
	546 => std_logic_vector(to_unsigned(42, 8)),
	547 => std_logic_vector(to_unsigned(42, 8)),
	548 => std_logic_vector(to_unsigned(41, 8)),
	549 => std_logic_vector(to_unsigned(42, 8)),
	550 => std_logic_vector(to_unsigned(42, 8)),
	551 => std_logic_vector(to_unsigned(41, 8)),
	552 => std_logic_vector(to_unsigned(42, 8)),
	553 => std_logic_vector(to_unsigned(42, 8)),
	554 => std_logic_vector(to_unsigned(41, 8)),
	555 => std_logic_vector(to_unsigned(42, 8)),
	556 => std_logic_vector(to_unsigned(42, 8)),
	557 => std_logic_vector(to_unsigned(41, 8)),
	558 => std_logic_vector(to_unsigned(42, 8)),
	559 => std_logic_vector(to_unsigned(42, 8)),
	560 => std_logic_vector(to_unsigned(42, 8)),
	561 => std_logic_vector(to_unsigned(42, 8)),
	562 => std_logic_vector(to_unsigned(42, 8)),
	563 => std_logic_vector(to_unsigned(41, 8)),
	564 => std_logic_vector(to_unsigned(41, 8)),
	565 => std_logic_vector(to_unsigned(41, 8)),
	566 => std_logic_vector(to_unsigned(42, 8)),
	567 => std_logic_vector(to_unsigned(42, 8)),
	568 => std_logic_vector(to_unsigned(42, 8)),
	569 => std_logic_vector(to_unsigned(41, 8)),
	570 => std_logic_vector(to_unsigned(42, 8)),
	571 => std_logic_vector(to_unsigned(41, 8)),
	572 => std_logic_vector(to_unsigned(41, 8)),
	573 => std_logic_vector(to_unsigned(42, 8)),
	574 => std_logic_vector(to_unsigned(41, 8)),
	575 => std_logic_vector(to_unsigned(42, 8)),
	576 => std_logic_vector(to_unsigned(42, 8)),
	577 => std_logic_vector(to_unsigned(41, 8)),
	578 => std_logic_vector(to_unsigned(41, 8)),
	579 => std_logic_vector(to_unsigned(41, 8)),
	580 => std_logic_vector(to_unsigned(41, 8)),
	581 => std_logic_vector(to_unsigned(42, 8)),
	582 => std_logic_vector(to_unsigned(42, 8)),
	583 => std_logic_vector(to_unsigned(42, 8)),
	584 => std_logic_vector(to_unsigned(41, 8)),
	585 => std_logic_vector(to_unsigned(42, 8)),
	586 => std_logic_vector(to_unsigned(41, 8)),
	587 => std_logic_vector(to_unsigned(41, 8)),
	588 => std_logic_vector(to_unsigned(41, 8)),
	589 => std_logic_vector(to_unsigned(42, 8)),
	590 => std_logic_vector(to_unsigned(41, 8)),
	591 => std_logic_vector(to_unsigned(41, 8)),
	592 => std_logic_vector(to_unsigned(41, 8)),
	593 => std_logic_vector(to_unsigned(41, 8)),
	594 => std_logic_vector(to_unsigned(41, 8)),
	595 => std_logic_vector(to_unsigned(42, 8)),
	596 => std_logic_vector(to_unsigned(41, 8)),
	597 => std_logic_vector(to_unsigned(41, 8)),
	598 => std_logic_vector(to_unsigned(41, 8)),
	599 => std_logic_vector(to_unsigned(41, 8)),
	600 => std_logic_vector(to_unsigned(42, 8)),
	601 => std_logic_vector(to_unsigned(42, 8)),
	602 => std_logic_vector(to_unsigned(42, 8)),
	603 => std_logic_vector(to_unsigned(42, 8)),
	604 => std_logic_vector(to_unsigned(42, 8)),
	605 => std_logic_vector(to_unsigned(41, 8)),
	606 => std_logic_vector(to_unsigned(41, 8)),
	607 => std_logic_vector(to_unsigned(42, 8)),
	608 => std_logic_vector(to_unsigned(42, 8)),
	609 => std_logic_vector(to_unsigned(41, 8)),
	610 => std_logic_vector(to_unsigned(41, 8)),
	611 => std_logic_vector(to_unsigned(42, 8)),
	612 => std_logic_vector(to_unsigned(41, 8)),
	613 => std_logic_vector(to_unsigned(42, 8)),
	614 => std_logic_vector(to_unsigned(42, 8)),
	615 => std_logic_vector(to_unsigned(42, 8)),
	616 => std_logic_vector(to_unsigned(42, 8)),
	617 => std_logic_vector(to_unsigned(41, 8)),
	618 => std_logic_vector(to_unsigned(41, 8)),
	619 => std_logic_vector(to_unsigned(42, 8)),
	620 => std_logic_vector(to_unsigned(41, 8)),
	621 => std_logic_vector(to_unsigned(42, 8)),
	622 => std_logic_vector(to_unsigned(41, 8)),
	623 => std_logic_vector(to_unsigned(41, 8)),
	624 => std_logic_vector(to_unsigned(42, 8)),
	625 => std_logic_vector(to_unsigned(42, 8)),
	626 => std_logic_vector(to_unsigned(42, 8)),
	627 => std_logic_vector(to_unsigned(42, 8)),
	628 => std_logic_vector(to_unsigned(41, 8)),
	629 => std_logic_vector(to_unsigned(41, 8)),
	630 => std_logic_vector(to_unsigned(42, 8)),
	631 => std_logic_vector(to_unsigned(42, 8)),
	632 => std_logic_vector(to_unsigned(42, 8)),
	633 => std_logic_vector(to_unsigned(42, 8)),
	634 => std_logic_vector(to_unsigned(41, 8)),
	635 => std_logic_vector(to_unsigned(41, 8)),
	636 => std_logic_vector(to_unsigned(41, 8)),
	637 => std_logic_vector(to_unsigned(42, 8)),
	638 => std_logic_vector(to_unsigned(42, 8)),
	639 => std_logic_vector(to_unsigned(41, 8)),
	640 => std_logic_vector(to_unsigned(41, 8)),
	641 => std_logic_vector(to_unsigned(41, 8)),
	642 => std_logic_vector(to_unsigned(42, 8)),
	643 => std_logic_vector(to_unsigned(42, 8)),
	644 => std_logic_vector(to_unsigned(42, 8)),
	645 => std_logic_vector(to_unsigned(41, 8)),
	646 => std_logic_vector(to_unsigned(42, 8)),
	647 => std_logic_vector(to_unsigned(41, 8)),
	648 => std_logic_vector(to_unsigned(42, 8)),
	649 => std_logic_vector(to_unsigned(42, 8)),
	650 => std_logic_vector(to_unsigned(41, 8)),
	651 => std_logic_vector(to_unsigned(42, 8)),
	652 => std_logic_vector(to_unsigned(41, 8)),
	653 => std_logic_vector(to_unsigned(41, 8)),
	654 => std_logic_vector(to_unsigned(41, 8)),
	655 => std_logic_vector(to_unsigned(41, 8)),
	656 => std_logic_vector(to_unsigned(42, 8)),
	657 => std_logic_vector(to_unsigned(42, 8)),
	658 => std_logic_vector(to_unsigned(42, 8)),
	659 => std_logic_vector(to_unsigned(41, 8)),
	660 => std_logic_vector(to_unsigned(41, 8)),
	661 => std_logic_vector(to_unsigned(42, 8)),
	662 => std_logic_vector(to_unsigned(41, 8)),
	663 => std_logic_vector(to_unsigned(41, 8)),
	664 => std_logic_vector(to_unsigned(41, 8)),
	665 => std_logic_vector(to_unsigned(42, 8)),
	666 => std_logic_vector(to_unsigned(42, 8)),
	667 => std_logic_vector(to_unsigned(42, 8)),
	668 => std_logic_vector(to_unsigned(42, 8)),
	669 => std_logic_vector(to_unsigned(41, 8)),
	670 => std_logic_vector(to_unsigned(41, 8)),
	671 => std_logic_vector(to_unsigned(41, 8)),
	672 => std_logic_vector(to_unsigned(41, 8)),
	673 => std_logic_vector(to_unsigned(42, 8)),
	674 => std_logic_vector(to_unsigned(41, 8)),
	675 => std_logic_vector(to_unsigned(42, 8)),
	676 => std_logic_vector(to_unsigned(41, 8)),
	677 => std_logic_vector(to_unsigned(41, 8)),
	678 => std_logic_vector(to_unsigned(42, 8)),
	679 => std_logic_vector(to_unsigned(41, 8)),
	680 => std_logic_vector(to_unsigned(42, 8)),
	681 => std_logic_vector(to_unsigned(41, 8)),
	682 => std_logic_vector(to_unsigned(42, 8)),
	683 => std_logic_vector(to_unsigned(41, 8)),
	684 => std_logic_vector(to_unsigned(42, 8)),
	685 => std_logic_vector(to_unsigned(42, 8)),
	686 => std_logic_vector(to_unsigned(42, 8)),
	687 => std_logic_vector(to_unsigned(41, 8)),
	688 => std_logic_vector(to_unsigned(42, 8)),
	689 => std_logic_vector(to_unsigned(41, 8)),
	690 => std_logic_vector(to_unsigned(41, 8)),
	691 => std_logic_vector(to_unsigned(41, 8)),
	692 => std_logic_vector(to_unsigned(41, 8)),
	693 => std_logic_vector(to_unsigned(41, 8)),
	694 => std_logic_vector(to_unsigned(42, 8)),
	695 => std_logic_vector(to_unsigned(42, 8)),
	696 => std_logic_vector(to_unsigned(41, 8)),
	697 => std_logic_vector(to_unsigned(42, 8)),
	698 => std_logic_vector(to_unsigned(42, 8)),
	699 => std_logic_vector(to_unsigned(41, 8)),
	700 => std_logic_vector(to_unsigned(42, 8)),
	701 => std_logic_vector(to_unsigned(41, 8)),
	702 => std_logic_vector(to_unsigned(41, 8)),
	703 => std_logic_vector(to_unsigned(41, 8)),
	704 => std_logic_vector(to_unsigned(42, 8)),
	705 => std_logic_vector(to_unsigned(41, 8)),
	706 => std_logic_vector(to_unsigned(41, 8)),
	707 => std_logic_vector(to_unsigned(41, 8)),
	708 => std_logic_vector(to_unsigned(42, 8)),
	709 => std_logic_vector(to_unsigned(42, 8)),
	710 => std_logic_vector(to_unsigned(42, 8)),
	711 => std_logic_vector(to_unsigned(41, 8)),
	712 => std_logic_vector(to_unsigned(42, 8)),
	713 => std_logic_vector(to_unsigned(42, 8)),
	714 => std_logic_vector(to_unsigned(42, 8)),
	715 => std_logic_vector(to_unsigned(41, 8)),
	716 => std_logic_vector(to_unsigned(41, 8)),
	717 => std_logic_vector(to_unsigned(41, 8)),
	718 => std_logic_vector(to_unsigned(42, 8)),
	719 => std_logic_vector(to_unsigned(42, 8)),
	720 => std_logic_vector(to_unsigned(42, 8)),
	721 => std_logic_vector(to_unsigned(42, 8)),
	722 => std_logic_vector(to_unsigned(42, 8)),
	723 => std_logic_vector(to_unsigned(41, 8)),
	724 => std_logic_vector(to_unsigned(42, 8)),
	725 => std_logic_vector(to_unsigned(41, 8)),
	726 => std_logic_vector(to_unsigned(42, 8)),
	727 => std_logic_vector(to_unsigned(42, 8)),
	728 => std_logic_vector(to_unsigned(42, 8)),
	729 => std_logic_vector(to_unsigned(42, 8)),
	730 => std_logic_vector(to_unsigned(41, 8)),
	731 => std_logic_vector(to_unsigned(42, 8)),
	732 => std_logic_vector(to_unsigned(42, 8)),
	733 => std_logic_vector(to_unsigned(42, 8)),
	734 => std_logic_vector(to_unsigned(41, 8)),
	735 => std_logic_vector(to_unsigned(41, 8)),
	736 => std_logic_vector(to_unsigned(42, 8)),
	737 => std_logic_vector(to_unsigned(42, 8)),
	738 => std_logic_vector(to_unsigned(42, 8)),
	739 => std_logic_vector(to_unsigned(41, 8)),
	740 => std_logic_vector(to_unsigned(42, 8)),
	741 => std_logic_vector(to_unsigned(42, 8)),
	742 => std_logic_vector(to_unsigned(41, 8)),
	743 => std_logic_vector(to_unsigned(42, 8)),
	744 => std_logic_vector(to_unsigned(42, 8)),
	745 => std_logic_vector(to_unsigned(41, 8)),
	746 => std_logic_vector(to_unsigned(41, 8)),
	747 => std_logic_vector(to_unsigned(41, 8)),
	748 => std_logic_vector(to_unsigned(42, 8)),
	749 => std_logic_vector(to_unsigned(42, 8)),
	750 => std_logic_vector(to_unsigned(41, 8)),
	751 => std_logic_vector(to_unsigned(41, 8)),
	752 => std_logic_vector(to_unsigned(41, 8)),
	753 => std_logic_vector(to_unsigned(41, 8)),
	754 => std_logic_vector(to_unsigned(41, 8)),
	755 => std_logic_vector(to_unsigned(41, 8)),
	756 => std_logic_vector(to_unsigned(42, 8)),
	757 => std_logic_vector(to_unsigned(42, 8)),
	758 => std_logic_vector(to_unsigned(41, 8)),
	759 => std_logic_vector(to_unsigned(41, 8)),
	760 => std_logic_vector(to_unsigned(41, 8)),
	761 => std_logic_vector(to_unsigned(41, 8)),
	762 => std_logic_vector(to_unsigned(41, 8)),
	763 => std_logic_vector(to_unsigned(41, 8)),
	764 => std_logic_vector(to_unsigned(42, 8)),
	765 => std_logic_vector(to_unsigned(41, 8)),
	766 => std_logic_vector(to_unsigned(42, 8)),
	767 => std_logic_vector(to_unsigned(42, 8)),
	768 => std_logic_vector(to_unsigned(41, 8)),
	769 => std_logic_vector(to_unsigned(41, 8)),
	770 => std_logic_vector(to_unsigned(41, 8)),
	771 => std_logic_vector(to_unsigned(41, 8)),
	772 => std_logic_vector(to_unsigned(42, 8)),
	773 => std_logic_vector(to_unsigned(42, 8)),
	774 => std_logic_vector(to_unsigned(41, 8)),
	775 => std_logic_vector(to_unsigned(41, 8)),
	776 => std_logic_vector(to_unsigned(41, 8)),
	777 => std_logic_vector(to_unsigned(41, 8)),
	778 => std_logic_vector(to_unsigned(41, 8)),
	779 => std_logic_vector(to_unsigned(41, 8)),
	780 => std_logic_vector(to_unsigned(41, 8)),
	781 => std_logic_vector(to_unsigned(42, 8)),
	782 => std_logic_vector(to_unsigned(41, 8)),
	783 => std_logic_vector(to_unsigned(42, 8)),
	784 => std_logic_vector(to_unsigned(42, 8)),
	785 => std_logic_vector(to_unsigned(41, 8)),
	786 => std_logic_vector(to_unsigned(42, 8)),
	787 => std_logic_vector(to_unsigned(41, 8)),
	788 => std_logic_vector(to_unsigned(42, 8)),
	789 => std_logic_vector(to_unsigned(42, 8)),
	790 => std_logic_vector(to_unsigned(42, 8)),
	791 => std_logic_vector(to_unsigned(41, 8)),
	792 => std_logic_vector(to_unsigned(42, 8)),
	793 => std_logic_vector(to_unsigned(41, 8)),
	794 => std_logic_vector(to_unsigned(41, 8)),
	795 => std_logic_vector(to_unsigned(42, 8)),
	796 => std_logic_vector(to_unsigned(42, 8)),
	797 => std_logic_vector(to_unsigned(42, 8)),
	798 => std_logic_vector(to_unsigned(41, 8)),
	799 => std_logic_vector(to_unsigned(42, 8)),
	800 => std_logic_vector(to_unsigned(42, 8)),
	801 => std_logic_vector(to_unsigned(41, 8)),
	802 => std_logic_vector(to_unsigned(42, 8)),
	803 => std_logic_vector(to_unsigned(41, 8)),
	804 => std_logic_vector(to_unsigned(41, 8)),
	805 => std_logic_vector(to_unsigned(41, 8)),
	806 => std_logic_vector(to_unsigned(41, 8)),
	807 => std_logic_vector(to_unsigned(41, 8)),
	808 => std_logic_vector(to_unsigned(41, 8)),
	809 => std_logic_vector(to_unsigned(42, 8)),
	810 => std_logic_vector(to_unsigned(42, 8)),
	811 => std_logic_vector(to_unsigned(42, 8)),
	812 => std_logic_vector(to_unsigned(41, 8)),
	813 => std_logic_vector(to_unsigned(41, 8)),
	814 => std_logic_vector(to_unsigned(42, 8)),
	815 => std_logic_vector(to_unsigned(41, 8)),
	816 => std_logic_vector(to_unsigned(42, 8)),
	817 => std_logic_vector(to_unsigned(42, 8)),
	818 => std_logic_vector(to_unsigned(42, 8)),
	819 => std_logic_vector(to_unsigned(41, 8)),
	820 => std_logic_vector(to_unsigned(42, 8)),
	821 => std_logic_vector(to_unsigned(42, 8)),
	822 => std_logic_vector(to_unsigned(41, 8)),
	823 => std_logic_vector(to_unsigned(41, 8)),
	824 => std_logic_vector(to_unsigned(42, 8)),
	825 => std_logic_vector(to_unsigned(41, 8)),
	826 => std_logic_vector(to_unsigned(41, 8)),
	827 => std_logic_vector(to_unsigned(41, 8)),
	828 => std_logic_vector(to_unsigned(42, 8)),
	829 => std_logic_vector(to_unsigned(42, 8)),
	830 => std_logic_vector(to_unsigned(42, 8)),
	831 => std_logic_vector(to_unsigned(42, 8)),
	832 => std_logic_vector(to_unsigned(41, 8)),
	833 => std_logic_vector(to_unsigned(41, 8)),
	834 => std_logic_vector(to_unsigned(42, 8)),
	835 => std_logic_vector(to_unsigned(41, 8)),
	836 => std_logic_vector(to_unsigned(42, 8)),
	837 => std_logic_vector(to_unsigned(42, 8)),
	838 => std_logic_vector(to_unsigned(42, 8)),
	839 => std_logic_vector(to_unsigned(42, 8)),
	840 => std_logic_vector(to_unsigned(42, 8)),
	841 => std_logic_vector(to_unsigned(41, 8)),
	842 => std_logic_vector(to_unsigned(41, 8)),
	843 => std_logic_vector(to_unsigned(42, 8)),
	844 => std_logic_vector(to_unsigned(41, 8)),
	845 => std_logic_vector(to_unsigned(41, 8)),
	846 => std_logic_vector(to_unsigned(41, 8)),
	847 => std_logic_vector(to_unsigned(42, 8)),
	848 => std_logic_vector(to_unsigned(42, 8)),
	849 => std_logic_vector(to_unsigned(42, 8)),
	850 => std_logic_vector(to_unsigned(42, 8)),
	851 => std_logic_vector(to_unsigned(41, 8)),
	852 => std_logic_vector(to_unsigned(41, 8)),
	853 => std_logic_vector(to_unsigned(41, 8)),
	854 => std_logic_vector(to_unsigned(41, 8)),
	855 => std_logic_vector(to_unsigned(42, 8)),
	856 => std_logic_vector(to_unsigned(42, 8)),
	857 => std_logic_vector(to_unsigned(42, 8)),
	858 => std_logic_vector(to_unsigned(41, 8)),
	859 => std_logic_vector(to_unsigned(41, 8)),
	860 => std_logic_vector(to_unsigned(42, 8)),
	861 => std_logic_vector(to_unsigned(42, 8)),
	862 => std_logic_vector(to_unsigned(42, 8)),
	863 => std_logic_vector(to_unsigned(41, 8)),
	864 => std_logic_vector(to_unsigned(42, 8)),
	865 => std_logic_vector(to_unsigned(42, 8)),
	866 => std_logic_vector(to_unsigned(41, 8)),
	867 => std_logic_vector(to_unsigned(41, 8)),
	868 => std_logic_vector(to_unsigned(41, 8)),
	869 => std_logic_vector(to_unsigned(42, 8)),
	870 => std_logic_vector(to_unsigned(42, 8)),
	871 => std_logic_vector(to_unsigned(42, 8)),
	872 => std_logic_vector(to_unsigned(41, 8)),
	873 => std_logic_vector(to_unsigned(42, 8)),
	874 => std_logic_vector(to_unsigned(42, 8)),
	875 => std_logic_vector(to_unsigned(41, 8)),
	876 => std_logic_vector(to_unsigned(41, 8)),
	877 => std_logic_vector(to_unsigned(42, 8)),
	878 => std_logic_vector(to_unsigned(42, 8)),
	879 => std_logic_vector(to_unsigned(41, 8)),
	880 => std_logic_vector(to_unsigned(41, 8)),
	881 => std_logic_vector(to_unsigned(42, 8)),
	882 => std_logic_vector(to_unsigned(42, 8)),
	883 => std_logic_vector(to_unsigned(41, 8)),
	884 => std_logic_vector(to_unsigned(42, 8)),
	885 => std_logic_vector(to_unsigned(41, 8)),
	886 => std_logic_vector(to_unsigned(42, 8)),
	887 => std_logic_vector(to_unsigned(41, 8)),
	888 => std_logic_vector(to_unsigned(42, 8)),
	889 => std_logic_vector(to_unsigned(41, 8)),
	890 => std_logic_vector(to_unsigned(41, 8)),
	891 => std_logic_vector(to_unsigned(42, 8)),
	892 => std_logic_vector(to_unsigned(41, 8)),
	893 => std_logic_vector(to_unsigned(41, 8)),
	894 => std_logic_vector(to_unsigned(41, 8)),
	895 => std_logic_vector(to_unsigned(41, 8)),
	896 => std_logic_vector(to_unsigned(42, 8)),
	897 => std_logic_vector(to_unsigned(41, 8)),
	898 => std_logic_vector(to_unsigned(42, 8)),
	899 => std_logic_vector(to_unsigned(41, 8)),
	900 => std_logic_vector(to_unsigned(41, 8)),
	901 => std_logic_vector(to_unsigned(42, 8)),
	902 => std_logic_vector(to_unsigned(41, 8)),
	903 => std_logic_vector(to_unsigned(41, 8)),
	904 => std_logic_vector(to_unsigned(41, 8)),
	905 => std_logic_vector(to_unsigned(41, 8)),
	906 => std_logic_vector(to_unsigned(42, 8)),
	907 => std_logic_vector(to_unsigned(42, 8)),
	908 => std_logic_vector(to_unsigned(42, 8)),
	909 => std_logic_vector(to_unsigned(41, 8)),
	910 => std_logic_vector(to_unsigned(41, 8)),
	911 => std_logic_vector(to_unsigned(41, 8)),
	912 => std_logic_vector(to_unsigned(42, 8)),
	913 => std_logic_vector(to_unsigned(41, 8)),
	914 => std_logic_vector(to_unsigned(42, 8)),
	915 => std_logic_vector(to_unsigned(42, 8)),
	916 => std_logic_vector(to_unsigned(41, 8)),
	917 => std_logic_vector(to_unsigned(41, 8)),
	918 => std_logic_vector(to_unsigned(42, 8)),
	919 => std_logic_vector(to_unsigned(42, 8)),
	920 => std_logic_vector(to_unsigned(42, 8)),
	921 => std_logic_vector(to_unsigned(42, 8)),
	922 => std_logic_vector(to_unsigned(41, 8)),
	923 => std_logic_vector(to_unsigned(41, 8)),
	924 => std_logic_vector(to_unsigned(41, 8)),
	925 => std_logic_vector(to_unsigned(41, 8)),
	926 => std_logic_vector(to_unsigned(41, 8)),
	927 => std_logic_vector(to_unsigned(42, 8)),
	928 => std_logic_vector(to_unsigned(42, 8)),
	929 => std_logic_vector(to_unsigned(41, 8)),
	930 => std_logic_vector(to_unsigned(42, 8)),
	931 => std_logic_vector(to_unsigned(41, 8)),
	932 => std_logic_vector(to_unsigned(42, 8)),
	933 => std_logic_vector(to_unsigned(42, 8)),
	934 => std_logic_vector(to_unsigned(41, 8)),
	935 => std_logic_vector(to_unsigned(41, 8)),
	936 => std_logic_vector(to_unsigned(42, 8)),
	937 => std_logic_vector(to_unsigned(41, 8)),
	938 => std_logic_vector(to_unsigned(41, 8)),
	939 => std_logic_vector(to_unsigned(42, 8)),
	940 => std_logic_vector(to_unsigned(42, 8)),
	941 => std_logic_vector(to_unsigned(42, 8)),
	942 => std_logic_vector(to_unsigned(41, 8)),
	943 => std_logic_vector(to_unsigned(41, 8)),
	944 => std_logic_vector(to_unsigned(41, 8)),
	945 => std_logic_vector(to_unsigned(42, 8)),
	946 => std_logic_vector(to_unsigned(41, 8)),
	947 => std_logic_vector(to_unsigned(42, 8)),
	948 => std_logic_vector(to_unsigned(41, 8)),
	949 => std_logic_vector(to_unsigned(41, 8)),
	950 => std_logic_vector(to_unsigned(42, 8)),
	951 => std_logic_vector(to_unsigned(42, 8)),
	952 => std_logic_vector(to_unsigned(42, 8)),
	953 => std_logic_vector(to_unsigned(42, 8)),
	954 => std_logic_vector(to_unsigned(42, 8)),
	955 => std_logic_vector(to_unsigned(41, 8)),
	956 => std_logic_vector(to_unsigned(41, 8)),
	957 => std_logic_vector(to_unsigned(41, 8)),
	958 => std_logic_vector(to_unsigned(42, 8)),
	959 => std_logic_vector(to_unsigned(42, 8)),
	960 => std_logic_vector(to_unsigned(41, 8)),
	961 => std_logic_vector(to_unsigned(41, 8)),
	962 => std_logic_vector(to_unsigned(41, 8)),
	963 => std_logic_vector(to_unsigned(42, 8)),
	964 => std_logic_vector(to_unsigned(42, 8)),
	965 => std_logic_vector(to_unsigned(41, 8)),
	966 => std_logic_vector(to_unsigned(42, 8)),
	967 => std_logic_vector(to_unsigned(42, 8)),
	968 => std_logic_vector(to_unsigned(42, 8)),
	969 => std_logic_vector(to_unsigned(41, 8)),
	970 => std_logic_vector(to_unsigned(41, 8)),
	971 => std_logic_vector(to_unsigned(42, 8)),
	972 => std_logic_vector(to_unsigned(42, 8)),
	973 => std_logic_vector(to_unsigned(41, 8)),
	974 => std_logic_vector(to_unsigned(42, 8)),
	975 => std_logic_vector(to_unsigned(41, 8)),
	976 => std_logic_vector(to_unsigned(42, 8)),
	977 => std_logic_vector(to_unsigned(41, 8)),
	978 => std_logic_vector(to_unsigned(42, 8)),
	979 => std_logic_vector(to_unsigned(41, 8)),
	980 => std_logic_vector(to_unsigned(41, 8)),
	981 => std_logic_vector(to_unsigned(41, 8)),
	982 => std_logic_vector(to_unsigned(41, 8)),
	983 => std_logic_vector(to_unsigned(41, 8)),
	984 => std_logic_vector(to_unsigned(41, 8)),
	985 => std_logic_vector(to_unsigned(41, 8)),
	986 => std_logic_vector(to_unsigned(42, 8)),
	987 => std_logic_vector(to_unsigned(42, 8)),
	988 => std_logic_vector(to_unsigned(42, 8)),
	989 => std_logic_vector(to_unsigned(41, 8)),
	990 => std_logic_vector(to_unsigned(42, 8)),
	991 => std_logic_vector(to_unsigned(41, 8)),
	992 => std_logic_vector(to_unsigned(42, 8)),
	993 => std_logic_vector(to_unsigned(41, 8)),
	994 => std_logic_vector(to_unsigned(41, 8)),
	995 => std_logic_vector(to_unsigned(41, 8)),
	996 => std_logic_vector(to_unsigned(41, 8)),
	997 => std_logic_vector(to_unsigned(42, 8)),
	998 => std_logic_vector(to_unsigned(42, 8)),
	999 => std_logic_vector(to_unsigned(42, 8)),
	1000 => std_logic_vector(to_unsigned(41, 8)),
	1001 => std_logic_vector(to_unsigned(42, 8)),
	1002 => std_logic_vector(to_unsigned(41, 8)),
	1003 => std_logic_vector(to_unsigned(41, 8)),
	1004 => std_logic_vector(to_unsigned(41, 8)),
	1005 => std_logic_vector(to_unsigned(41, 8)),
	1006 => std_logic_vector(to_unsigned(42, 8)),
	1007 => std_logic_vector(to_unsigned(41, 8)),
	1008 => std_logic_vector(to_unsigned(41, 8)),
	1009 => std_logic_vector(to_unsigned(41, 8)),
	1010 => std_logic_vector(to_unsigned(42, 8)),
	1011 => std_logic_vector(to_unsigned(41, 8)),
	1012 => std_logic_vector(to_unsigned(42, 8)),
	1013 => std_logic_vector(to_unsigned(42, 8)),
	1014 => std_logic_vector(to_unsigned(42, 8)),
	1015 => std_logic_vector(to_unsigned(42, 8)),
	1016 => std_logic_vector(to_unsigned(41, 8)),
	1017 => std_logic_vector(to_unsigned(42, 8)),
	1018 => std_logic_vector(to_unsigned(42, 8)),
	1019 => std_logic_vector(to_unsigned(41, 8)),
	1020 => std_logic_vector(to_unsigned(42, 8)),
	1021 => std_logic_vector(to_unsigned(41, 8)),
	1022 => std_logic_vector(to_unsigned(41, 8)),
	1023 => std_logic_vector(to_unsigned(41, 8)),
	1024 => std_logic_vector(to_unsigned(42, 8)),
	1025 => std_logic_vector(to_unsigned(42, 8)),
	1026 => std_logic_vector(to_unsigned(41, 8)),
	1027 => std_logic_vector(to_unsigned(42, 8)),
	1028 => std_logic_vector(to_unsigned(41, 8)),
	1029 => std_logic_vector(to_unsigned(42, 8)),
	1030 => std_logic_vector(to_unsigned(41, 8)),
	1031 => std_logic_vector(to_unsigned(42, 8)),
	1032 => std_logic_vector(to_unsigned(42, 8)),
	1033 => std_logic_vector(to_unsigned(42, 8)),
	1034 => std_logic_vector(to_unsigned(42, 8)),
	1035 => std_logic_vector(to_unsigned(41, 8)),
	1036 => std_logic_vector(to_unsigned(41, 8)),
	1037 => std_logic_vector(to_unsigned(41, 8)),
	1038 => std_logic_vector(to_unsigned(41, 8)),
	1039 => std_logic_vector(to_unsigned(41, 8)),
	1040 => std_logic_vector(to_unsigned(41, 8)),
	1041 => std_logic_vector(to_unsigned(41, 8)),
	1042 => std_logic_vector(to_unsigned(41, 8)),
	1043 => std_logic_vector(to_unsigned(41, 8)),
	1044 => std_logic_vector(to_unsigned(42, 8)),
	1045 => std_logic_vector(to_unsigned(41, 8)),
	1046 => std_logic_vector(to_unsigned(41, 8)),
	1047 => std_logic_vector(to_unsigned(41, 8)),
	1048 => std_logic_vector(to_unsigned(41, 8)),
	1049 => std_logic_vector(to_unsigned(41, 8)),
	1050 => std_logic_vector(to_unsigned(41, 8)),
	1051 => std_logic_vector(to_unsigned(41, 8)),
	1052 => std_logic_vector(to_unsigned(41, 8)),
	1053 => std_logic_vector(to_unsigned(41, 8)),
	1054 => std_logic_vector(to_unsigned(42, 8)),
	1055 => std_logic_vector(to_unsigned(42, 8)),
	1056 => std_logic_vector(to_unsigned(41, 8)),
	1057 => std_logic_vector(to_unsigned(41, 8)),
	1058 => std_logic_vector(to_unsigned(41, 8)),
	1059 => std_logic_vector(to_unsigned(41, 8)),
	1060 => std_logic_vector(to_unsigned(42, 8)),
	1061 => std_logic_vector(to_unsigned(41, 8)),
	1062 => std_logic_vector(to_unsigned(41, 8)),
	1063 => std_logic_vector(to_unsigned(41, 8)),
	1064 => std_logic_vector(to_unsigned(41, 8)),
	1065 => std_logic_vector(to_unsigned(41, 8)),
	1066 => std_logic_vector(to_unsigned(41, 8)),
	1067 => std_logic_vector(to_unsigned(42, 8)),
	1068 => std_logic_vector(to_unsigned(42, 8)),
	1069 => std_logic_vector(to_unsigned(42, 8)),
	1070 => std_logic_vector(to_unsigned(41, 8)),
	1071 => std_logic_vector(to_unsigned(41, 8)),
	1072 => std_logic_vector(to_unsigned(42, 8)),
	1073 => std_logic_vector(to_unsigned(41, 8)),
	1074 => std_logic_vector(to_unsigned(41, 8)),
	1075 => std_logic_vector(to_unsigned(42, 8)),
	1076 => std_logic_vector(to_unsigned(41, 8)),
	1077 => std_logic_vector(to_unsigned(41, 8)),
	1078 => std_logic_vector(to_unsigned(41, 8)),
	1079 => std_logic_vector(to_unsigned(41, 8)),
	1080 => std_logic_vector(to_unsigned(42, 8)),
	1081 => std_logic_vector(to_unsigned(41, 8)),
	1082 => std_logic_vector(to_unsigned(42, 8)),
	1083 => std_logic_vector(to_unsigned(42, 8)),
	1084 => std_logic_vector(to_unsigned(41, 8)),
	1085 => std_logic_vector(to_unsigned(41, 8)),
	1086 => std_logic_vector(to_unsigned(42, 8)),
	1087 => std_logic_vector(to_unsigned(41, 8)),
	1088 => std_logic_vector(to_unsigned(41, 8)),
	1089 => std_logic_vector(to_unsigned(41, 8)),
	1090 => std_logic_vector(to_unsigned(42, 8)),
	1091 => std_logic_vector(to_unsigned(41, 8)),
	1092 => std_logic_vector(to_unsigned(42, 8)),
	1093 => std_logic_vector(to_unsigned(41, 8)),
	1094 => std_logic_vector(to_unsigned(41, 8)),
	1095 => std_logic_vector(to_unsigned(42, 8)),
	1096 => std_logic_vector(to_unsigned(41, 8)),
	1097 => std_logic_vector(to_unsigned(41, 8)),
	1098 => std_logic_vector(to_unsigned(41, 8)),
	1099 => std_logic_vector(to_unsigned(42, 8)),
	1100 => std_logic_vector(to_unsigned(41, 8)),
	1101 => std_logic_vector(to_unsigned(41, 8)),
	1102 => std_logic_vector(to_unsigned(42, 8)),
	1103 => std_logic_vector(to_unsigned(42, 8)),
	1104 => std_logic_vector(to_unsigned(41, 8)),
	1105 => std_logic_vector(to_unsigned(42, 8)),
	1106 => std_logic_vector(to_unsigned(42, 8)),
	1107 => std_logic_vector(to_unsigned(42, 8)),
	1108 => std_logic_vector(to_unsigned(41, 8)),
	1109 => std_logic_vector(to_unsigned(41, 8)),
	1110 => std_logic_vector(to_unsigned(42, 8)),
	1111 => std_logic_vector(to_unsigned(41, 8)),
	1112 => std_logic_vector(to_unsigned(42, 8)),
	1113 => std_logic_vector(to_unsigned(42, 8)),
	1114 => std_logic_vector(to_unsigned(41, 8)),
	1115 => std_logic_vector(to_unsigned(41, 8)),
	1116 => std_logic_vector(to_unsigned(42, 8)),
	1117 => std_logic_vector(to_unsigned(42, 8)),
	1118 => std_logic_vector(to_unsigned(41, 8)),
	1119 => std_logic_vector(to_unsigned(41, 8)),
	1120 => std_logic_vector(to_unsigned(41, 8)),
	1121 => std_logic_vector(to_unsigned(42, 8)),
	1122 => std_logic_vector(to_unsigned(41, 8)),
	1123 => std_logic_vector(to_unsigned(41, 8)),
	1124 => std_logic_vector(to_unsigned(42, 8)),
	1125 => std_logic_vector(to_unsigned(41, 8)),
	1126 => std_logic_vector(to_unsigned(42, 8)),
	1127 => std_logic_vector(to_unsigned(42, 8)),
	1128 => std_logic_vector(to_unsigned(41, 8)),
	1129 => std_logic_vector(to_unsigned(42, 8)),
	1130 => std_logic_vector(to_unsigned(41, 8)),
	1131 => std_logic_vector(to_unsigned(42, 8)),
	1132 => std_logic_vector(to_unsigned(42, 8)),
	1133 => std_logic_vector(to_unsigned(42, 8)),
	1134 => std_logic_vector(to_unsigned(42, 8)),
	1135 => std_logic_vector(to_unsigned(41, 8)),
	1136 => std_logic_vector(to_unsigned(42, 8)),
	1137 => std_logic_vector(to_unsigned(41, 8)),
	1138 => std_logic_vector(to_unsigned(41, 8)),
	1139 => std_logic_vector(to_unsigned(41, 8)),
	1140 => std_logic_vector(to_unsigned(41, 8)),
	1141 => std_logic_vector(to_unsigned(41, 8)),
	1142 => std_logic_vector(to_unsigned(41, 8)),
	1143 => std_logic_vector(to_unsigned(41, 8)),
	1144 => std_logic_vector(to_unsigned(42, 8)),
	1145 => std_logic_vector(to_unsigned(42, 8)),
	1146 => std_logic_vector(to_unsigned(41, 8)),
	1147 => std_logic_vector(to_unsigned(41, 8)),
	1148 => std_logic_vector(to_unsigned(41, 8)),
	1149 => std_logic_vector(to_unsigned(41, 8)),
	1150 => std_logic_vector(to_unsigned(41, 8)),
	1151 => std_logic_vector(to_unsigned(41, 8)),
	1152 => std_logic_vector(to_unsigned(42, 8)),
	1153 => std_logic_vector(to_unsigned(42, 8)),
	1154 => std_logic_vector(to_unsigned(41, 8)),
	1155 => std_logic_vector(to_unsigned(42, 8)),
	1156 => std_logic_vector(to_unsigned(42, 8)),
	1157 => std_logic_vector(to_unsigned(42, 8)),
	1158 => std_logic_vector(to_unsigned(42, 8)),
	1159 => std_logic_vector(to_unsigned(42, 8)),
	1160 => std_logic_vector(to_unsigned(41, 8)),
	1161 => std_logic_vector(to_unsigned(41, 8)),
	1162 => std_logic_vector(to_unsigned(41, 8)),
	1163 => std_logic_vector(to_unsigned(41, 8)),
	1164 => std_logic_vector(to_unsigned(42, 8)),
	1165 => std_logic_vector(to_unsigned(41, 8)),
	1166 => std_logic_vector(to_unsigned(42, 8)),
	1167 => std_logic_vector(to_unsigned(41, 8)),
	1168 => std_logic_vector(to_unsigned(42, 8)),
	1169 => std_logic_vector(to_unsigned(42, 8)),
	1170 => std_logic_vector(to_unsigned(42, 8)),
	1171 => std_logic_vector(to_unsigned(41, 8)),
	1172 => std_logic_vector(to_unsigned(41, 8)),
	1173 => std_logic_vector(to_unsigned(42, 8)),
	1174 => std_logic_vector(to_unsigned(41, 8)),
	1175 => std_logic_vector(to_unsigned(42, 8)),
	1176 => std_logic_vector(to_unsigned(42, 8)),
	1177 => std_logic_vector(to_unsigned(42, 8)),
	1178 => std_logic_vector(to_unsigned(41, 8)),
	1179 => std_logic_vector(to_unsigned(42, 8)),
	1180 => std_logic_vector(to_unsigned(41, 8)),
	1181 => std_logic_vector(to_unsigned(42, 8)),
	1182 => std_logic_vector(to_unsigned(42, 8)),
	1183 => std_logic_vector(to_unsigned(41, 8)),
	1184 => std_logic_vector(to_unsigned(42, 8)),
	1185 => std_logic_vector(to_unsigned(41, 8)),
	1186 => std_logic_vector(to_unsigned(41, 8)),
	1187 => std_logic_vector(to_unsigned(42, 8)),
	1188 => std_logic_vector(to_unsigned(42, 8)),
	1189 => std_logic_vector(to_unsigned(41, 8)),
	1190 => std_logic_vector(to_unsigned(42, 8)),
	1191 => std_logic_vector(to_unsigned(41, 8)),
	1192 => std_logic_vector(to_unsigned(41, 8)),
	1193 => std_logic_vector(to_unsigned(41, 8)),
	1194 => std_logic_vector(to_unsigned(42, 8)),
	1195 => std_logic_vector(to_unsigned(41, 8)),
	1196 => std_logic_vector(to_unsigned(42, 8)),
	1197 => std_logic_vector(to_unsigned(42, 8)),
	1198 => std_logic_vector(to_unsigned(41, 8)),
	1199 => std_logic_vector(to_unsigned(42, 8)),
	1200 => std_logic_vector(to_unsigned(41, 8)),
	1201 => std_logic_vector(to_unsigned(41, 8)),
	1202 => std_logic_vector(to_unsigned(41, 8)),
	1203 => std_logic_vector(to_unsigned(42, 8)),
	1204 => std_logic_vector(to_unsigned(41, 8)),
	1205 => std_logic_vector(to_unsigned(42, 8)),
	1206 => std_logic_vector(to_unsigned(41, 8)),
	1207 => std_logic_vector(to_unsigned(42, 8)),
	1208 => std_logic_vector(to_unsigned(42, 8)),
	1209 => std_logic_vector(to_unsigned(41, 8)),
	1210 => std_logic_vector(to_unsigned(42, 8)),
	1211 => std_logic_vector(to_unsigned(41, 8)),
	1212 => std_logic_vector(to_unsigned(41, 8)),
	1213 => std_logic_vector(to_unsigned(42, 8)),
	1214 => std_logic_vector(to_unsigned(41, 8)),
	1215 => std_logic_vector(to_unsigned(41, 8)),
	1216 => std_logic_vector(to_unsigned(42, 8)),
	1217 => std_logic_vector(to_unsigned(41, 8)),
	1218 => std_logic_vector(to_unsigned(41, 8)),
	1219 => std_logic_vector(to_unsigned(42, 8)),
	1220 => std_logic_vector(to_unsigned(42, 8)),
	1221 => std_logic_vector(to_unsigned(41, 8)),
	1222 => std_logic_vector(to_unsigned(42, 8)),
	1223 => std_logic_vector(to_unsigned(41, 8)),
	1224 => std_logic_vector(to_unsigned(41, 8)),
	1225 => std_logic_vector(to_unsigned(41, 8)),
	1226 => std_logic_vector(to_unsigned(41, 8)),
	1227 => std_logic_vector(to_unsigned(42, 8)),
	1228 => std_logic_vector(to_unsigned(41, 8)),
	1229 => std_logic_vector(to_unsigned(42, 8)),
	1230 => std_logic_vector(to_unsigned(41, 8)),
	1231 => std_logic_vector(to_unsigned(41, 8)),
	1232 => std_logic_vector(to_unsigned(42, 8)),
	1233 => std_logic_vector(to_unsigned(41, 8)),
	1234 => std_logic_vector(to_unsigned(41, 8)),
	1235 => std_logic_vector(to_unsigned(42, 8)),
	1236 => std_logic_vector(to_unsigned(42, 8)),
	1237 => std_logic_vector(to_unsigned(41, 8)),
	1238 => std_logic_vector(to_unsigned(41, 8)),
	1239 => std_logic_vector(to_unsigned(42, 8)),
	1240 => std_logic_vector(to_unsigned(42, 8)),
	1241 => std_logic_vector(to_unsigned(42, 8)),
	1242 => std_logic_vector(to_unsigned(42, 8)),
	1243 => std_logic_vector(to_unsigned(42, 8)),
	1244 => std_logic_vector(to_unsigned(42, 8)),
	1245 => std_logic_vector(to_unsigned(42, 8)),
	1246 => std_logic_vector(to_unsigned(41, 8)),
	1247 => std_logic_vector(to_unsigned(41, 8)),
	1248 => std_logic_vector(to_unsigned(42, 8)),
	1249 => std_logic_vector(to_unsigned(42, 8)),
	1250 => std_logic_vector(to_unsigned(42, 8)),
	1251 => std_logic_vector(to_unsigned(42, 8)),
	1252 => std_logic_vector(to_unsigned(42, 8)),
	1253 => std_logic_vector(to_unsigned(41, 8)),
	1254 => std_logic_vector(to_unsigned(42, 8)),
	1255 => std_logic_vector(to_unsigned(41, 8)),
	1256 => std_logic_vector(to_unsigned(41, 8)),
	1257 => std_logic_vector(to_unsigned(42, 8)),
	1258 => std_logic_vector(to_unsigned(41, 8)),
	1259 => std_logic_vector(to_unsigned(41, 8)),
	1260 => std_logic_vector(to_unsigned(42, 8)),
	1261 => std_logic_vector(to_unsigned(42, 8)),
	1262 => std_logic_vector(to_unsigned(42, 8)),
	1263 => std_logic_vector(to_unsigned(41, 8)),
	1264 => std_logic_vector(to_unsigned(41, 8)),
	1265 => std_logic_vector(to_unsigned(42, 8)),
	1266 => std_logic_vector(to_unsigned(41, 8)),
	1267 => std_logic_vector(to_unsigned(42, 8)),
	1268 => std_logic_vector(to_unsigned(42, 8)),
	1269 => std_logic_vector(to_unsigned(41, 8)),
	1270 => std_logic_vector(to_unsigned(42, 8)),
	1271 => std_logic_vector(to_unsigned(41, 8)),
	1272 => std_logic_vector(to_unsigned(42, 8)),
	1273 => std_logic_vector(to_unsigned(41, 8)),
	1274 => std_logic_vector(to_unsigned(42, 8)),
	1275 => std_logic_vector(to_unsigned(41, 8)),
	1276 => std_logic_vector(to_unsigned(42, 8)),
	1277 => std_logic_vector(to_unsigned(41, 8)),
	1278 => std_logic_vector(to_unsigned(41, 8)),
	1279 => std_logic_vector(to_unsigned(42, 8)),
	1280 => std_logic_vector(to_unsigned(41, 8)),
	1281 => std_logic_vector(to_unsigned(41, 8)),
	1282 => std_logic_vector(to_unsigned(41, 8)),
	1283 => std_logic_vector(to_unsigned(42, 8)),
	1284 => std_logic_vector(to_unsigned(41, 8)),
	1285 => std_logic_vector(to_unsigned(42, 8)),
	1286 => std_logic_vector(to_unsigned(42, 8)),
	1287 => std_logic_vector(to_unsigned(42, 8)),
	1288 => std_logic_vector(to_unsigned(41, 8)),
	1289 => std_logic_vector(to_unsigned(41, 8)),
	1290 => std_logic_vector(to_unsigned(41, 8)),
	1291 => std_logic_vector(to_unsigned(42, 8)),
	1292 => std_logic_vector(to_unsigned(41, 8)),
	1293 => std_logic_vector(to_unsigned(42, 8)),
	1294 => std_logic_vector(to_unsigned(42, 8)),
	1295 => std_logic_vector(to_unsigned(42, 8)),
	1296 => std_logic_vector(to_unsigned(42, 8)),
	1297 => std_logic_vector(to_unsigned(42, 8)),
	1298 => std_logic_vector(to_unsigned(41, 8)),
	1299 => std_logic_vector(to_unsigned(41, 8)),
	1300 => std_logic_vector(to_unsigned(42, 8)),
	1301 => std_logic_vector(to_unsigned(42, 8)),
	1302 => std_logic_vector(to_unsigned(42, 8)),
	1303 => std_logic_vector(to_unsigned(41, 8)),
	1304 => std_logic_vector(to_unsigned(41, 8)),
	1305 => std_logic_vector(to_unsigned(41, 8)),
	1306 => std_logic_vector(to_unsigned(42, 8)),
	1307 => std_logic_vector(to_unsigned(41, 8)),
	1308 => std_logic_vector(to_unsigned(41, 8)),
	1309 => std_logic_vector(to_unsigned(42, 8)),
	1310 => std_logic_vector(to_unsigned(42, 8)),
	1311 => std_logic_vector(to_unsigned(42, 8)),
	1312 => std_logic_vector(to_unsigned(42, 8)),
	1313 => std_logic_vector(to_unsigned(41, 8)),
	1314 => std_logic_vector(to_unsigned(41, 8)),
	1315 => std_logic_vector(to_unsigned(42, 8)),
	1316 => std_logic_vector(to_unsigned(42, 8)),
	1317 => std_logic_vector(to_unsigned(42, 8)),
	1318 => std_logic_vector(to_unsigned(42, 8)),
	1319 => std_logic_vector(to_unsigned(42, 8)),
	1320 => std_logic_vector(to_unsigned(41, 8)),
	1321 => std_logic_vector(to_unsigned(42, 8)),
	1322 => std_logic_vector(to_unsigned(42, 8)),
	1323 => std_logic_vector(to_unsigned(41, 8)),
	1324 => std_logic_vector(to_unsigned(42, 8)),
	1325 => std_logic_vector(to_unsigned(41, 8)),
	1326 => std_logic_vector(to_unsigned(42, 8)),
	1327 => std_logic_vector(to_unsigned(41, 8)),
	1328 => std_logic_vector(to_unsigned(41, 8)),
	1329 => std_logic_vector(to_unsigned(42, 8)),
	1330 => std_logic_vector(to_unsigned(42, 8)),
	1331 => std_logic_vector(to_unsigned(41, 8)),
	1332 => std_logic_vector(to_unsigned(42, 8)),
	1333 => std_logic_vector(to_unsigned(41, 8)),
	1334 => std_logic_vector(to_unsigned(42, 8)),
	1335 => std_logic_vector(to_unsigned(42, 8)),
	1336 => std_logic_vector(to_unsigned(42, 8)),
	1337 => std_logic_vector(to_unsigned(42, 8)),
	1338 => std_logic_vector(to_unsigned(41, 8)),
	1339 => std_logic_vector(to_unsigned(42, 8)),
	1340 => std_logic_vector(to_unsigned(41, 8)),
	1341 => std_logic_vector(to_unsigned(41, 8)),
	1342 => std_logic_vector(to_unsigned(41, 8)),
	1343 => std_logic_vector(to_unsigned(42, 8)),
	1344 => std_logic_vector(to_unsigned(41, 8)),
	1345 => std_logic_vector(to_unsigned(41, 8)),
	1346 => std_logic_vector(to_unsigned(42, 8)),
	1347 => std_logic_vector(to_unsigned(42, 8)),
	1348 => std_logic_vector(to_unsigned(41, 8)),
	1349 => std_logic_vector(to_unsigned(41, 8)),
	1350 => std_logic_vector(to_unsigned(42, 8)),
	1351 => std_logic_vector(to_unsigned(42, 8)),
	1352 => std_logic_vector(to_unsigned(42, 8)),
	1353 => std_logic_vector(to_unsigned(41, 8)),
	1354 => std_logic_vector(to_unsigned(41, 8)),
	1355 => std_logic_vector(to_unsigned(42, 8)),
	1356 => std_logic_vector(to_unsigned(41, 8)),
	1357 => std_logic_vector(to_unsigned(42, 8)),
	1358 => std_logic_vector(to_unsigned(42, 8)),
	1359 => std_logic_vector(to_unsigned(41, 8)),
	1360 => std_logic_vector(to_unsigned(42, 8)),
	1361 => std_logic_vector(to_unsigned(42, 8)),
	1362 => std_logic_vector(to_unsigned(42, 8)),
	1363 => std_logic_vector(to_unsigned(41, 8)),
	1364 => std_logic_vector(to_unsigned(41, 8)),
	1365 => std_logic_vector(to_unsigned(42, 8)),
	1366 => std_logic_vector(to_unsigned(42, 8)),
	1367 => std_logic_vector(to_unsigned(42, 8)),
	1368 => std_logic_vector(to_unsigned(41, 8)),
	1369 => std_logic_vector(to_unsigned(42, 8)),
	1370 => std_logic_vector(to_unsigned(42, 8)),
	1371 => std_logic_vector(to_unsigned(41, 8)),
	1372 => std_logic_vector(to_unsigned(41, 8)),
	1373 => std_logic_vector(to_unsigned(41, 8)),
	1374 => std_logic_vector(to_unsigned(42, 8)),
	1375 => std_logic_vector(to_unsigned(41, 8)),
	1376 => std_logic_vector(to_unsigned(42, 8)),
	1377 => std_logic_vector(to_unsigned(42, 8)),
	1378 => std_logic_vector(to_unsigned(42, 8)),
	1379 => std_logic_vector(to_unsigned(42, 8)),
	1380 => std_logic_vector(to_unsigned(42, 8)),
	1381 => std_logic_vector(to_unsigned(41, 8)),
	1382 => std_logic_vector(to_unsigned(42, 8)),
	1383 => std_logic_vector(to_unsigned(41, 8)),
	1384 => std_logic_vector(to_unsigned(41, 8)),
	1385 => std_logic_vector(to_unsigned(42, 8)),
	1386 => std_logic_vector(to_unsigned(41, 8)),
	1387 => std_logic_vector(to_unsigned(42, 8)),
	1388 => std_logic_vector(to_unsigned(42, 8)),
	1389 => std_logic_vector(to_unsigned(41, 8)),
	1390 => std_logic_vector(to_unsigned(41, 8)),
	1391 => std_logic_vector(to_unsigned(42, 8)),
	1392 => std_logic_vector(to_unsigned(41, 8)),
	1393 => std_logic_vector(to_unsigned(41, 8)),
	1394 => std_logic_vector(to_unsigned(42, 8)),
	1395 => std_logic_vector(to_unsigned(41, 8)),
	1396 => std_logic_vector(to_unsigned(42, 8)),
	1397 => std_logic_vector(to_unsigned(41, 8)),
	1398 => std_logic_vector(to_unsigned(41, 8)),
	1399 => std_logic_vector(to_unsigned(42, 8)),
	1400 => std_logic_vector(to_unsigned(41, 8)),
	1401 => std_logic_vector(to_unsigned(41, 8)),
	1402 => std_logic_vector(to_unsigned(42, 8)),
	1403 => std_logic_vector(to_unsigned(42, 8)),
	1404 => std_logic_vector(to_unsigned(41, 8)),
	1405 => std_logic_vector(to_unsigned(41, 8)),
	1406 => std_logic_vector(to_unsigned(42, 8)),
	1407 => std_logic_vector(to_unsigned(42, 8)),
	1408 => std_logic_vector(to_unsigned(42, 8)),
	1409 => std_logic_vector(to_unsigned(41, 8)),
	1410 => std_logic_vector(to_unsigned(42, 8)),
	1411 => std_logic_vector(to_unsigned(41, 8)),
	1412 => std_logic_vector(to_unsigned(42, 8)),
	1413 => std_logic_vector(to_unsigned(42, 8)),
	1414 => std_logic_vector(to_unsigned(42, 8)),
	1415 => std_logic_vector(to_unsigned(42, 8)),
	1416 => std_logic_vector(to_unsigned(41, 8)),
	1417 => std_logic_vector(to_unsigned(41, 8)),
	1418 => std_logic_vector(to_unsigned(42, 8)),
	1419 => std_logic_vector(to_unsigned(42, 8)),
	1420 => std_logic_vector(to_unsigned(42, 8)),
	1421 => std_logic_vector(to_unsigned(42, 8)),
	1422 => std_logic_vector(to_unsigned(41, 8)),
	1423 => std_logic_vector(to_unsigned(41, 8)),
	1424 => std_logic_vector(to_unsigned(42, 8)),
	1425 => std_logic_vector(to_unsigned(41, 8)),
	1426 => std_logic_vector(to_unsigned(42, 8)),
	1427 => std_logic_vector(to_unsigned(42, 8)),
	1428 => std_logic_vector(to_unsigned(41, 8)),
	1429 => std_logic_vector(to_unsigned(41, 8)),
	1430 => std_logic_vector(to_unsigned(42, 8)),
	1431 => std_logic_vector(to_unsigned(41, 8)),
	1432 => std_logic_vector(to_unsigned(41, 8)),
	1433 => std_logic_vector(to_unsigned(42, 8)),
	1434 => std_logic_vector(to_unsigned(41, 8)),
	1435 => std_logic_vector(to_unsigned(41, 8)),
	1436 => std_logic_vector(to_unsigned(42, 8)),
	1437 => std_logic_vector(to_unsigned(41, 8)),
	1438 => std_logic_vector(to_unsigned(41, 8)),
	1439 => std_logic_vector(to_unsigned(42, 8)),
	1440 => std_logic_vector(to_unsigned(42, 8)),
	1441 => std_logic_vector(to_unsigned(42, 8)),
	1442 => std_logic_vector(to_unsigned(41, 8)),
	1443 => std_logic_vector(to_unsigned(42, 8)),
	1444 => std_logic_vector(to_unsigned(41, 8)),
	1445 => std_logic_vector(to_unsigned(41, 8)),
	1446 => std_logic_vector(to_unsigned(41, 8)),
	1447 => std_logic_vector(to_unsigned(41, 8)),
	1448 => std_logic_vector(to_unsigned(42, 8)),
	1449 => std_logic_vector(to_unsigned(42, 8)),
	1450 => std_logic_vector(to_unsigned(41, 8)),
	1451 => std_logic_vector(to_unsigned(41, 8)),
	1452 => std_logic_vector(to_unsigned(42, 8)),
	1453 => std_logic_vector(to_unsigned(42, 8)),
	1454 => std_logic_vector(to_unsigned(41, 8)),
	1455 => std_logic_vector(to_unsigned(41, 8)),
	1456 => std_logic_vector(to_unsigned(42, 8)),
	1457 => std_logic_vector(to_unsigned(42, 8)),
	1458 => std_logic_vector(to_unsigned(41, 8)),
	1459 => std_logic_vector(to_unsigned(42, 8)),
	1460 => std_logic_vector(to_unsigned(42, 8)),
	1461 => std_logic_vector(to_unsigned(41, 8)),
	1462 => std_logic_vector(to_unsigned(41, 8)),
	1463 => std_logic_vector(to_unsigned(41, 8)),
	1464 => std_logic_vector(to_unsigned(41, 8)),
	1465 => std_logic_vector(to_unsigned(41, 8)),
	1466 => std_logic_vector(to_unsigned(42, 8)),
	1467 => std_logic_vector(to_unsigned(41, 8)),
	1468 => std_logic_vector(to_unsigned(41, 8)),
	1469 => std_logic_vector(to_unsigned(42, 8)),
	1470 => std_logic_vector(to_unsigned(41, 8)),
	1471 => std_logic_vector(to_unsigned(41, 8)),
	1472 => std_logic_vector(to_unsigned(42, 8)),
	1473 => std_logic_vector(to_unsigned(42, 8)),
	1474 => std_logic_vector(to_unsigned(41, 8)),
	1475 => std_logic_vector(to_unsigned(42, 8)),
	1476 => std_logic_vector(to_unsigned(41, 8)),
	1477 => std_logic_vector(to_unsigned(42, 8)),
	1478 => std_logic_vector(to_unsigned(42, 8)),
	1479 => std_logic_vector(to_unsigned(41, 8)),
	1480 => std_logic_vector(to_unsigned(41, 8)),
	1481 => std_logic_vector(to_unsigned(42, 8)),
	1482 => std_logic_vector(to_unsigned(42, 8)),
	1483 => std_logic_vector(to_unsigned(42, 8)),
	1484 => std_logic_vector(to_unsigned(41, 8)),
	1485 => std_logic_vector(to_unsigned(42, 8)),
	1486 => std_logic_vector(to_unsigned(41, 8)),
	1487 => std_logic_vector(to_unsigned(41, 8)),
	1488 => std_logic_vector(to_unsigned(41, 8)),
	1489 => std_logic_vector(to_unsigned(41, 8)),
	1490 => std_logic_vector(to_unsigned(42, 8)),
	1491 => std_logic_vector(to_unsigned(41, 8)),
	1492 => std_logic_vector(to_unsigned(41, 8)),
	1493 => std_logic_vector(to_unsigned(41, 8)),
	1494 => std_logic_vector(to_unsigned(41, 8)),
	1495 => std_logic_vector(to_unsigned(42, 8)),
	1496 => std_logic_vector(to_unsigned(41, 8)),
	1497 => std_logic_vector(to_unsigned(41, 8)),
	1498 => std_logic_vector(to_unsigned(42, 8)),
	1499 => std_logic_vector(to_unsigned(41, 8)),
	1500 => std_logic_vector(to_unsigned(41, 8)),
	1501 => std_logic_vector(to_unsigned(41, 8)),
	1502 => std_logic_vector(to_unsigned(41, 8)),
	1503 => std_logic_vector(to_unsigned(42, 8)),
	1504 => std_logic_vector(to_unsigned(41, 8)),
	1505 => std_logic_vector(to_unsigned(42, 8)),
	1506 => std_logic_vector(to_unsigned(42, 8)),
	1507 => std_logic_vector(to_unsigned(42, 8)),
	1508 => std_logic_vector(to_unsigned(41, 8)),
	1509 => std_logic_vector(to_unsigned(41, 8)),
	1510 => std_logic_vector(to_unsigned(41, 8)),
	1511 => std_logic_vector(to_unsigned(42, 8)),
	1512 => std_logic_vector(to_unsigned(42, 8)),
	1513 => std_logic_vector(to_unsigned(41, 8)),
	1514 => std_logic_vector(to_unsigned(42, 8)),
	1515 => std_logic_vector(to_unsigned(42, 8)),
	1516 => std_logic_vector(to_unsigned(41, 8)),
	1517 => std_logic_vector(to_unsigned(42, 8)),
	1518 => std_logic_vector(to_unsigned(42, 8)),
	1519 => std_logic_vector(to_unsigned(41, 8)),
	1520 => std_logic_vector(to_unsigned(41, 8)),
	1521 => std_logic_vector(to_unsigned(41, 8)),
	1522 => std_logic_vector(to_unsigned(42, 8)),
	1523 => std_logic_vector(to_unsigned(42, 8)),
	1524 => std_logic_vector(to_unsigned(41, 8)),
	1525 => std_logic_vector(to_unsigned(42, 8)),
	1526 => std_logic_vector(to_unsigned(42, 8)),
	1527 => std_logic_vector(to_unsigned(42, 8)),
	1528 => std_logic_vector(to_unsigned(41, 8)),
	1529 => std_logic_vector(to_unsigned(42, 8)),
	1530 => std_logic_vector(to_unsigned(42, 8)),
	1531 => std_logic_vector(to_unsigned(41, 8)),
	1532 => std_logic_vector(to_unsigned(41, 8)),
	1533 => std_logic_vector(to_unsigned(41, 8)),
	1534 => std_logic_vector(to_unsigned(42, 8)),
	1535 => std_logic_vector(to_unsigned(41, 8)),
	1536 => std_logic_vector(to_unsigned(41, 8)),
	1537 => std_logic_vector(to_unsigned(41, 8)),
	1538 => std_logic_vector(to_unsigned(41, 8)),
	1539 => std_logic_vector(to_unsigned(41, 8)),
	1540 => std_logic_vector(to_unsigned(42, 8)),
	1541 => std_logic_vector(to_unsigned(41, 8)),
	1542 => std_logic_vector(to_unsigned(41, 8)),
	1543 => std_logic_vector(to_unsigned(41, 8)),
	1544 => std_logic_vector(to_unsigned(41, 8)),
	1545 => std_logic_vector(to_unsigned(42, 8)),
	1546 => std_logic_vector(to_unsigned(41, 8)),
	1547 => std_logic_vector(to_unsigned(42, 8)),
	1548 => std_logic_vector(to_unsigned(42, 8)),
	1549 => std_logic_vector(to_unsigned(42, 8)),
	1550 => std_logic_vector(to_unsigned(42, 8)),
	1551 => std_logic_vector(to_unsigned(41, 8)),
	1552 => std_logic_vector(to_unsigned(41, 8)),
	1553 => std_logic_vector(to_unsigned(41, 8)),
	1554 => std_logic_vector(to_unsigned(42, 8)),
	1555 => std_logic_vector(to_unsigned(42, 8)),
	1556 => std_logic_vector(to_unsigned(42, 8)),
	1557 => std_logic_vector(to_unsigned(42, 8)),
	1558 => std_logic_vector(to_unsigned(41, 8)),
	1559 => std_logic_vector(to_unsigned(42, 8)),
	1560 => std_logic_vector(to_unsigned(42, 8)),
	1561 => std_logic_vector(to_unsigned(41, 8)),
	1562 => std_logic_vector(to_unsigned(42, 8)),
	1563 => std_logic_vector(to_unsigned(42, 8)),
	1564 => std_logic_vector(to_unsigned(41, 8)),
	1565 => std_logic_vector(to_unsigned(42, 8)),
	1566 => std_logic_vector(to_unsigned(41, 8)),
	1567 => std_logic_vector(to_unsigned(41, 8)),
	1568 => std_logic_vector(to_unsigned(42, 8)),
	1569 => std_logic_vector(to_unsigned(41, 8)),
	1570 => std_logic_vector(to_unsigned(42, 8)),
	1571 => std_logic_vector(to_unsigned(42, 8)),
	1572 => std_logic_vector(to_unsigned(42, 8)),
	1573 => std_logic_vector(to_unsigned(41, 8)),
	1574 => std_logic_vector(to_unsigned(42, 8)),
	1575 => std_logic_vector(to_unsigned(42, 8)),
	1576 => std_logic_vector(to_unsigned(41, 8)),
	1577 => std_logic_vector(to_unsigned(42, 8)),
	1578 => std_logic_vector(to_unsigned(41, 8)),
	1579 => std_logic_vector(to_unsigned(42, 8)),
	1580 => std_logic_vector(to_unsigned(41, 8)),
	1581 => std_logic_vector(to_unsigned(41, 8)),
	1582 => std_logic_vector(to_unsigned(42, 8)),
	1583 => std_logic_vector(to_unsigned(42, 8)),
	1584 => std_logic_vector(to_unsigned(41, 8)),
	1585 => std_logic_vector(to_unsigned(41, 8)),
	1586 => std_logic_vector(to_unsigned(41, 8)),
	1587 => std_logic_vector(to_unsigned(41, 8)),
	1588 => std_logic_vector(to_unsigned(42, 8)),
	1589 => std_logic_vector(to_unsigned(42, 8)),
	1590 => std_logic_vector(to_unsigned(42, 8)),
	1591 => std_logic_vector(to_unsigned(41, 8)),
	1592 => std_logic_vector(to_unsigned(41, 8)),
	1593 => std_logic_vector(to_unsigned(42, 8)),
	1594 => std_logic_vector(to_unsigned(42, 8)),
	1595 => std_logic_vector(to_unsigned(42, 8)),
	1596 => std_logic_vector(to_unsigned(42, 8)),
	1597 => std_logic_vector(to_unsigned(41, 8)),
	1598 => std_logic_vector(to_unsigned(41, 8)),
	1599 => std_logic_vector(to_unsigned(42, 8)),
	1600 => std_logic_vector(to_unsigned(41, 8)),
	1601 => std_logic_vector(to_unsigned(42, 8)),
	1602 => std_logic_vector(to_unsigned(42, 8)),
	1603 => std_logic_vector(to_unsigned(42, 8)),
	1604 => std_logic_vector(to_unsigned(42, 8)),
	1605 => std_logic_vector(to_unsigned(41, 8)),
	1606 => std_logic_vector(to_unsigned(42, 8)),
	1607 => std_logic_vector(to_unsigned(42, 8)),
	1608 => std_logic_vector(to_unsigned(42, 8)),
	1609 => std_logic_vector(to_unsigned(42, 8)),
	1610 => std_logic_vector(to_unsigned(41, 8)),
	1611 => std_logic_vector(to_unsigned(42, 8)),
	1612 => std_logic_vector(to_unsigned(41, 8)),
	1613 => std_logic_vector(to_unsigned(41, 8)),
	1614 => std_logic_vector(to_unsigned(42, 8)),
	1615 => std_logic_vector(to_unsigned(42, 8)),
	1616 => std_logic_vector(to_unsigned(42, 8)),
	1617 => std_logic_vector(to_unsigned(41, 8)),
	1618 => std_logic_vector(to_unsigned(41, 8)),
	1619 => std_logic_vector(to_unsigned(42, 8)),
	1620 => std_logic_vector(to_unsigned(42, 8)),
	1621 => std_logic_vector(to_unsigned(42, 8)),
	1622 => std_logic_vector(to_unsigned(41, 8)),
	1623 => std_logic_vector(to_unsigned(42, 8)),
	1624 => std_logic_vector(to_unsigned(41, 8)),
	1625 => std_logic_vector(to_unsigned(41, 8)),
	1626 => std_logic_vector(to_unsigned(42, 8)),
	1627 => std_logic_vector(to_unsigned(41, 8)),
	1628 => std_logic_vector(to_unsigned(42, 8)),
	1629 => std_logic_vector(to_unsigned(41, 8)),
	1630 => std_logic_vector(to_unsigned(42, 8)),
	1631 => std_logic_vector(to_unsigned(42, 8)),
	1632 => std_logic_vector(to_unsigned(42, 8)),
	1633 => std_logic_vector(to_unsigned(42, 8)),
	1634 => std_logic_vector(to_unsigned(42, 8)),
	1635 => std_logic_vector(to_unsigned(42, 8)),
	1636 => std_logic_vector(to_unsigned(41, 8)),
	1637 => std_logic_vector(to_unsigned(41, 8)),
	1638 => std_logic_vector(to_unsigned(42, 8)),
	1639 => std_logic_vector(to_unsigned(41, 8)),
	1640 => std_logic_vector(to_unsigned(41, 8)),
	1641 => std_logic_vector(to_unsigned(42, 8)),
	1642 => std_logic_vector(to_unsigned(41, 8)),
	1643 => std_logic_vector(to_unsigned(41, 8)),
	1644 => std_logic_vector(to_unsigned(42, 8)),
	1645 => std_logic_vector(to_unsigned(42, 8)),
	1646 => std_logic_vector(to_unsigned(42, 8)),
	1647 => std_logic_vector(to_unsigned(42, 8)),
	1648 => std_logic_vector(to_unsigned(41, 8)),
	1649 => std_logic_vector(to_unsigned(41, 8)),
	1650 => std_logic_vector(to_unsigned(42, 8)),
	1651 => std_logic_vector(to_unsigned(41, 8)),
	1652 => std_logic_vector(to_unsigned(42, 8)),
	1653 => std_logic_vector(to_unsigned(42, 8)),
	1654 => std_logic_vector(to_unsigned(42, 8)),
	1655 => std_logic_vector(to_unsigned(41, 8)),
	1656 => std_logic_vector(to_unsigned(41, 8)),
	1657 => std_logic_vector(to_unsigned(42, 8)),
	1658 => std_logic_vector(to_unsigned(42, 8)),
	1659 => std_logic_vector(to_unsigned(41, 8)),
	1660 => std_logic_vector(to_unsigned(42, 8)),
	1661 => std_logic_vector(to_unsigned(41, 8)),
	1662 => std_logic_vector(to_unsigned(41, 8)),
	1663 => std_logic_vector(to_unsigned(42, 8)),
	1664 => std_logic_vector(to_unsigned(41, 8)),
	1665 => std_logic_vector(to_unsigned(41, 8)),
	1666 => std_logic_vector(to_unsigned(41, 8)),
	1667 => std_logic_vector(to_unsigned(41, 8)),
	1668 => std_logic_vector(to_unsigned(41, 8)),
	1669 => std_logic_vector(to_unsigned(41, 8)),
	1670 => std_logic_vector(to_unsigned(42, 8)),
	1671 => std_logic_vector(to_unsigned(42, 8)),
	1672 => std_logic_vector(to_unsigned(42, 8)),
	1673 => std_logic_vector(to_unsigned(42, 8)),
	1674 => std_logic_vector(to_unsigned(41, 8)),
	1675 => std_logic_vector(to_unsigned(42, 8)),
	1676 => std_logic_vector(to_unsigned(41, 8)),
	1677 => std_logic_vector(to_unsigned(42, 8)),
	1678 => std_logic_vector(to_unsigned(42, 8)),
	1679 => std_logic_vector(to_unsigned(42, 8)),
	1680 => std_logic_vector(to_unsigned(41, 8)),
	1681 => std_logic_vector(to_unsigned(41, 8)),
	1682 => std_logic_vector(to_unsigned(42, 8)),
	1683 => std_logic_vector(to_unsigned(42, 8)),
	1684 => std_logic_vector(to_unsigned(41, 8)),
	1685 => std_logic_vector(to_unsigned(42, 8)),
	1686 => std_logic_vector(to_unsigned(42, 8)),
	1687 => std_logic_vector(to_unsigned(41, 8)),
	1688 => std_logic_vector(to_unsigned(42, 8)),
	1689 => std_logic_vector(to_unsigned(42, 8)),
	1690 => std_logic_vector(to_unsigned(41, 8)),
	1691 => std_logic_vector(to_unsigned(41, 8)),
	1692 => std_logic_vector(to_unsigned(41, 8)),
	1693 => std_logic_vector(to_unsigned(41, 8)),
	1694 => std_logic_vector(to_unsigned(41, 8)),
	1695 => std_logic_vector(to_unsigned(42, 8)),
	1696 => std_logic_vector(to_unsigned(41, 8)),
	1697 => std_logic_vector(to_unsigned(42, 8)),
	1698 => std_logic_vector(to_unsigned(42, 8)),
	1699 => std_logic_vector(to_unsigned(41, 8)),
	1700 => std_logic_vector(to_unsigned(42, 8)),
	1701 => std_logic_vector(to_unsigned(41, 8)),
	1702 => std_logic_vector(to_unsigned(42, 8)),
	1703 => std_logic_vector(to_unsigned(42, 8)),
	1704 => std_logic_vector(to_unsigned(42, 8)),
	1705 => std_logic_vector(to_unsigned(42, 8)),
	1706 => std_logic_vector(to_unsigned(42, 8)),
	1707 => std_logic_vector(to_unsigned(42, 8)),
	1708 => std_logic_vector(to_unsigned(42, 8)),
	1709 => std_logic_vector(to_unsigned(41, 8)),
	1710 => std_logic_vector(to_unsigned(41, 8)),
	1711 => std_logic_vector(to_unsigned(41, 8)),
	1712 => std_logic_vector(to_unsigned(41, 8)),
	1713 => std_logic_vector(to_unsigned(41, 8)),
	1714 => std_logic_vector(to_unsigned(41, 8)),
	1715 => std_logic_vector(to_unsigned(41, 8)),
	1716 => std_logic_vector(to_unsigned(41, 8)),
	1717 => std_logic_vector(to_unsigned(41, 8)),
	1718 => std_logic_vector(to_unsigned(41, 8)),
	1719 => std_logic_vector(to_unsigned(41, 8)),
	1720 => std_logic_vector(to_unsigned(41, 8)),
	1721 => std_logic_vector(to_unsigned(41, 8)),
	1722 => std_logic_vector(to_unsigned(42, 8)),
	1723 => std_logic_vector(to_unsigned(42, 8)),
	1724 => std_logic_vector(to_unsigned(42, 8)),
	1725 => std_logic_vector(to_unsigned(41, 8)),
	1726 => std_logic_vector(to_unsigned(41, 8)),
	1727 => std_logic_vector(to_unsigned(41, 8)),
	1728 => std_logic_vector(to_unsigned(42, 8)),
	1729 => std_logic_vector(to_unsigned(41, 8)),
	1730 => std_logic_vector(to_unsigned(42, 8)),
	1731 => std_logic_vector(to_unsigned(41, 8)),
	1732 => std_logic_vector(to_unsigned(42, 8)),
	1733 => std_logic_vector(to_unsigned(41, 8)),
	1734 => std_logic_vector(to_unsigned(42, 8)),
	1735 => std_logic_vector(to_unsigned(41, 8)),
	1736 => std_logic_vector(to_unsigned(42, 8)),
	1737 => std_logic_vector(to_unsigned(41, 8)),
	1738 => std_logic_vector(to_unsigned(41, 8)),
	1739 => std_logic_vector(to_unsigned(41, 8)),
	1740 => std_logic_vector(to_unsigned(42, 8)),
	1741 => std_logic_vector(to_unsigned(41, 8)),
	1742 => std_logic_vector(to_unsigned(42, 8)),
	1743 => std_logic_vector(to_unsigned(41, 8)),
	1744 => std_logic_vector(to_unsigned(42, 8)),
	1745 => std_logic_vector(to_unsigned(41, 8)),
	1746 => std_logic_vector(to_unsigned(42, 8)),
	1747 => std_logic_vector(to_unsigned(42, 8)),
	1748 => std_logic_vector(to_unsigned(42, 8)),
	1749 => std_logic_vector(to_unsigned(41, 8)),
	1750 => std_logic_vector(to_unsigned(42, 8)),
	1751 => std_logic_vector(to_unsigned(42, 8)),
	1752 => std_logic_vector(to_unsigned(41, 8)),
	1753 => std_logic_vector(to_unsigned(41, 8)),
	1754 => std_logic_vector(to_unsigned(42, 8)),
	1755 => std_logic_vector(to_unsigned(42, 8)),
	1756 => std_logic_vector(to_unsigned(42, 8)),
	1757 => std_logic_vector(to_unsigned(41, 8)),
	1758 => std_logic_vector(to_unsigned(41, 8)),
	1759 => std_logic_vector(to_unsigned(42, 8)),
	1760 => std_logic_vector(to_unsigned(41, 8)),
	1761 => std_logic_vector(to_unsigned(41, 8)),
	1762 => std_logic_vector(to_unsigned(41, 8)),
	1763 => std_logic_vector(to_unsigned(42, 8)),
	1764 => std_logic_vector(to_unsigned(41, 8)),
	1765 => std_logic_vector(to_unsigned(42, 8)),
	1766 => std_logic_vector(to_unsigned(42, 8)),
	1767 => std_logic_vector(to_unsigned(42, 8)),
	1768 => std_logic_vector(to_unsigned(42, 8)),
	1769 => std_logic_vector(to_unsigned(41, 8)),
	1770 => std_logic_vector(to_unsigned(41, 8)),
	1771 => std_logic_vector(to_unsigned(41, 8)),
	1772 => std_logic_vector(to_unsigned(41, 8)),
	1773 => std_logic_vector(to_unsigned(42, 8)),
	1774 => std_logic_vector(to_unsigned(42, 8)),
	1775 => std_logic_vector(to_unsigned(42, 8)),
	1776 => std_logic_vector(to_unsigned(41, 8)),
	1777 => std_logic_vector(to_unsigned(41, 8)),
	1778 => std_logic_vector(to_unsigned(42, 8)),
	1779 => std_logic_vector(to_unsigned(42, 8)),
	1780 => std_logic_vector(to_unsigned(42, 8)),
	1781 => std_logic_vector(to_unsigned(41, 8)),
	1782 => std_logic_vector(to_unsigned(42, 8)),
	1783 => std_logic_vector(to_unsigned(41, 8)),
	1784 => std_logic_vector(to_unsigned(42, 8)),
	1785 => std_logic_vector(to_unsigned(41, 8)),
	1786 => std_logic_vector(to_unsigned(42, 8)),
	1787 => std_logic_vector(to_unsigned(42, 8)),
	1788 => std_logic_vector(to_unsigned(41, 8)),
	1789 => std_logic_vector(to_unsigned(41, 8)),
	1790 => std_logic_vector(to_unsigned(42, 8)),
	1791 => std_logic_vector(to_unsigned(41, 8)),
	1792 => std_logic_vector(to_unsigned(41, 8)),
	1793 => std_logic_vector(to_unsigned(42, 8)),
	1794 => std_logic_vector(to_unsigned(42, 8)),
	1795 => std_logic_vector(to_unsigned(41, 8)),
	1796 => std_logic_vector(to_unsigned(41, 8)),
	1797 => std_logic_vector(to_unsigned(42, 8)),
	1798 => std_logic_vector(to_unsigned(42, 8)),
	1799 => std_logic_vector(to_unsigned(42, 8)),
	1800 => std_logic_vector(to_unsigned(42, 8)),
	1801 => std_logic_vector(to_unsigned(42, 8)),
	1802 => std_logic_vector(to_unsigned(42, 8)),
	1803 => std_logic_vector(to_unsigned(41, 8)),
	1804 => std_logic_vector(to_unsigned(42, 8)),
	1805 => std_logic_vector(to_unsigned(41, 8)),
	1806 => std_logic_vector(to_unsigned(42, 8)),
	1807 => std_logic_vector(to_unsigned(41, 8)),
	1808 => std_logic_vector(to_unsigned(42, 8)),
	1809 => std_logic_vector(to_unsigned(41, 8)),
	1810 => std_logic_vector(to_unsigned(41, 8)),
	1811 => std_logic_vector(to_unsigned(42, 8)),
	1812 => std_logic_vector(to_unsigned(42, 8)),
	1813 => std_logic_vector(to_unsigned(41, 8)),
	1814 => std_logic_vector(to_unsigned(42, 8)),
	1815 => std_logic_vector(to_unsigned(42, 8)),
	1816 => std_logic_vector(to_unsigned(42, 8)),
	1817 => std_logic_vector(to_unsigned(42, 8)),
	1818 => std_logic_vector(to_unsigned(41, 8)),
	1819 => std_logic_vector(to_unsigned(41, 8)),
	1820 => std_logic_vector(to_unsigned(42, 8)),
	1821 => std_logic_vector(to_unsigned(41, 8)),
	1822 => std_logic_vector(to_unsigned(41, 8)),
	1823 => std_logic_vector(to_unsigned(41, 8)),
	1824 => std_logic_vector(to_unsigned(41, 8)),
	1825 => std_logic_vector(to_unsigned(41, 8)),
	1826 => std_logic_vector(to_unsigned(42, 8)),
	1827 => std_logic_vector(to_unsigned(41, 8)),
	1828 => std_logic_vector(to_unsigned(42, 8)),
	1829 => std_logic_vector(to_unsigned(41, 8)),
	1830 => std_logic_vector(to_unsigned(41, 8)),
	1831 => std_logic_vector(to_unsigned(41, 8)),
	1832 => std_logic_vector(to_unsigned(41, 8)),
	1833 => std_logic_vector(to_unsigned(41, 8)),
	1834 => std_logic_vector(to_unsigned(41, 8)),
	1835 => std_logic_vector(to_unsigned(41, 8)),
	1836 => std_logic_vector(to_unsigned(41, 8)),
	1837 => std_logic_vector(to_unsigned(42, 8)),
	1838 => std_logic_vector(to_unsigned(42, 8)),
	1839 => std_logic_vector(to_unsigned(42, 8)),
	1840 => std_logic_vector(to_unsigned(41, 8)),
	1841 => std_logic_vector(to_unsigned(41, 8)),
	1842 => std_logic_vector(to_unsigned(42, 8)),
	1843 => std_logic_vector(to_unsigned(41, 8)),
	1844 => std_logic_vector(to_unsigned(41, 8)),
	1845 => std_logic_vector(to_unsigned(42, 8)),
	1846 => std_logic_vector(to_unsigned(42, 8)),
	1847 => std_logic_vector(to_unsigned(41, 8)),
	1848 => std_logic_vector(to_unsigned(41, 8)),
	1849 => std_logic_vector(to_unsigned(41, 8)),
	1850 => std_logic_vector(to_unsigned(41, 8)),
	1851 => std_logic_vector(to_unsigned(42, 8)),
	1852 => std_logic_vector(to_unsigned(42, 8)),
	1853 => std_logic_vector(to_unsigned(41, 8)),
	1854 => std_logic_vector(to_unsigned(42, 8)),
	1855 => std_logic_vector(to_unsigned(42, 8)),
	1856 => std_logic_vector(to_unsigned(42, 8)),
	1857 => std_logic_vector(to_unsigned(41, 8)),
	1858 => std_logic_vector(to_unsigned(41, 8)),
	1859 => std_logic_vector(to_unsigned(42, 8)),
	1860 => std_logic_vector(to_unsigned(42, 8)),
	1861 => std_logic_vector(to_unsigned(41, 8)),
	1862 => std_logic_vector(to_unsigned(42, 8)),
	1863 => std_logic_vector(to_unsigned(41, 8)),
	1864 => std_logic_vector(to_unsigned(41, 8)),
	1865 => std_logic_vector(to_unsigned(41, 8)),
	1866 => std_logic_vector(to_unsigned(42, 8)),
	1867 => std_logic_vector(to_unsigned(42, 8)),
	1868 => std_logic_vector(to_unsigned(41, 8)),
	1869 => std_logic_vector(to_unsigned(41, 8)),
	1870 => std_logic_vector(to_unsigned(42, 8)),
	1871 => std_logic_vector(to_unsigned(41, 8)),
	1872 => std_logic_vector(to_unsigned(41, 8)),
	1873 => std_logic_vector(to_unsigned(41, 8)),
	1874 => std_logic_vector(to_unsigned(41, 8)),
	1875 => std_logic_vector(to_unsigned(41, 8)),
	1876 => std_logic_vector(to_unsigned(42, 8)),
	1877 => std_logic_vector(to_unsigned(41, 8)),
	1878 => std_logic_vector(to_unsigned(42, 8)),
	1879 => std_logic_vector(to_unsigned(42, 8)),
	1880 => std_logic_vector(to_unsigned(41, 8)),
	1881 => std_logic_vector(to_unsigned(42, 8)),
	1882 => std_logic_vector(to_unsigned(41, 8)),
	1883 => std_logic_vector(to_unsigned(42, 8)),
	1884 => std_logic_vector(to_unsigned(42, 8)),
	1885 => std_logic_vector(to_unsigned(41, 8)),
	1886 => std_logic_vector(to_unsigned(42, 8)),
	1887 => std_logic_vector(to_unsigned(42, 8)),
	1888 => std_logic_vector(to_unsigned(42, 8)),
	1889 => std_logic_vector(to_unsigned(42, 8)),
	1890 => std_logic_vector(to_unsigned(42, 8)),
	1891 => std_logic_vector(to_unsigned(42, 8)),
	1892 => std_logic_vector(to_unsigned(41, 8)),
	1893 => std_logic_vector(to_unsigned(42, 8)),
	1894 => std_logic_vector(to_unsigned(41, 8)),
	1895 => std_logic_vector(to_unsigned(41, 8)),
	1896 => std_logic_vector(to_unsigned(42, 8)),
	1897 => std_logic_vector(to_unsigned(41, 8)),
	1898 => std_logic_vector(to_unsigned(41, 8)),
	1899 => std_logic_vector(to_unsigned(42, 8)),
	1900 => std_logic_vector(to_unsigned(42, 8)),
	1901 => std_logic_vector(to_unsigned(42, 8)),
	1902 => std_logic_vector(to_unsigned(42, 8)),
	1903 => std_logic_vector(to_unsigned(41, 8)),
	1904 => std_logic_vector(to_unsigned(42, 8)),
	1905 => std_logic_vector(to_unsigned(42, 8)),
	1906 => std_logic_vector(to_unsigned(41, 8)),
	1907 => std_logic_vector(to_unsigned(41, 8)),
	1908 => std_logic_vector(to_unsigned(42, 8)),
	1909 => std_logic_vector(to_unsigned(41, 8)),
	1910 => std_logic_vector(to_unsigned(41, 8)),
	1911 => std_logic_vector(to_unsigned(41, 8)),
	1912 => std_logic_vector(to_unsigned(42, 8)),
	1913 => std_logic_vector(to_unsigned(42, 8)),
	1914 => std_logic_vector(to_unsigned(42, 8)),
	1915 => std_logic_vector(to_unsigned(42, 8)),
	1916 => std_logic_vector(to_unsigned(42, 8)),
	1917 => std_logic_vector(to_unsigned(41, 8)),
	1918 => std_logic_vector(to_unsigned(42, 8)),
	1919 => std_logic_vector(to_unsigned(41, 8)),
	1920 => std_logic_vector(to_unsigned(41, 8)),
	1921 => std_logic_vector(to_unsigned(41, 8)),
	1922 => std_logic_vector(to_unsigned(41, 8)),
	1923 => std_logic_vector(to_unsigned(42, 8)),
	1924 => std_logic_vector(to_unsigned(41, 8)),
	1925 => std_logic_vector(to_unsigned(41, 8)),
	1926 => std_logic_vector(to_unsigned(41, 8)),
	1927 => std_logic_vector(to_unsigned(42, 8)),
	1928 => std_logic_vector(to_unsigned(42, 8)),
	1929 => std_logic_vector(to_unsigned(42, 8)),
	1930 => std_logic_vector(to_unsigned(41, 8)),
	1931 => std_logic_vector(to_unsigned(41, 8)),
	1932 => std_logic_vector(to_unsigned(41, 8)),
	1933 => std_logic_vector(to_unsigned(42, 8)),
	1934 => std_logic_vector(to_unsigned(42, 8)),
	1935 => std_logic_vector(to_unsigned(41, 8)),
	1936 => std_logic_vector(to_unsigned(42, 8)),
	1937 => std_logic_vector(to_unsigned(41, 8)),
	1938 => std_logic_vector(to_unsigned(41, 8)),
	1939 => std_logic_vector(to_unsigned(42, 8)),
	1940 => std_logic_vector(to_unsigned(41, 8)),
	1941 => std_logic_vector(to_unsigned(42, 8)),
	1942 => std_logic_vector(to_unsigned(41, 8)),
	1943 => std_logic_vector(to_unsigned(41, 8)),
	1944 => std_logic_vector(to_unsigned(42, 8)),
	1945 => std_logic_vector(to_unsigned(42, 8)),
	1946 => std_logic_vector(to_unsigned(42, 8)),
	1947 => std_logic_vector(to_unsigned(41, 8)),
	1948 => std_logic_vector(to_unsigned(41, 8)),
	1949 => std_logic_vector(to_unsigned(41, 8)),
	1950 => std_logic_vector(to_unsigned(42, 8)),
	1951 => std_logic_vector(to_unsigned(42, 8)),
	1952 => std_logic_vector(to_unsigned(41, 8)),
	1953 => std_logic_vector(to_unsigned(41, 8)),
	1954 => std_logic_vector(to_unsigned(42, 8)),
	1955 => std_logic_vector(to_unsigned(42, 8)),
	1956 => std_logic_vector(to_unsigned(42, 8)),
	1957 => std_logic_vector(to_unsigned(42, 8)),
	1958 => std_logic_vector(to_unsigned(41, 8)),
	1959 => std_logic_vector(to_unsigned(41, 8)),
	1960 => std_logic_vector(to_unsigned(41, 8)),
	1961 => std_logic_vector(to_unsigned(42, 8)),
	1962 => std_logic_vector(to_unsigned(42, 8)),
	1963 => std_logic_vector(to_unsigned(41, 8)),
	1964 => std_logic_vector(to_unsigned(41, 8)),
	1965 => std_logic_vector(to_unsigned(42, 8)),
	1966 => std_logic_vector(to_unsigned(41, 8)),
	1967 => std_logic_vector(to_unsigned(41, 8)),
	1968 => std_logic_vector(to_unsigned(41, 8)),
	1969 => std_logic_vector(to_unsigned(41, 8)),
	1970 => std_logic_vector(to_unsigned(42, 8)),
	1971 => std_logic_vector(to_unsigned(42, 8)),
	1972 => std_logic_vector(to_unsigned(41, 8)),
	1973 => std_logic_vector(to_unsigned(41, 8)),
	1974 => std_logic_vector(to_unsigned(41, 8)),
	1975 => std_logic_vector(to_unsigned(42, 8)),
	1976 => std_logic_vector(to_unsigned(41, 8)),
	1977 => std_logic_vector(to_unsigned(41, 8)),
	1978 => std_logic_vector(to_unsigned(42, 8)),
	1979 => std_logic_vector(to_unsigned(41, 8)),
	1980 => std_logic_vector(to_unsigned(42, 8)),
	1981 => std_logic_vector(to_unsigned(41, 8)),
	1982 => std_logic_vector(to_unsigned(42, 8)),
	1983 => std_logic_vector(to_unsigned(41, 8)),
	1984 => std_logic_vector(to_unsigned(42, 8)),
	1985 => std_logic_vector(to_unsigned(41, 8)),
	1986 => std_logic_vector(to_unsigned(42, 8)),
	1987 => std_logic_vector(to_unsigned(42, 8)),
	1988 => std_logic_vector(to_unsigned(41, 8)),
	1989 => std_logic_vector(to_unsigned(42, 8)),
	1990 => std_logic_vector(to_unsigned(42, 8)),
	1991 => std_logic_vector(to_unsigned(42, 8)),
	1992 => std_logic_vector(to_unsigned(42, 8)),
	1993 => std_logic_vector(to_unsigned(41, 8)),
	1994 => std_logic_vector(to_unsigned(41, 8)),
	1995 => std_logic_vector(to_unsigned(42, 8)),
	1996 => std_logic_vector(to_unsigned(42, 8)),
	1997 => std_logic_vector(to_unsigned(42, 8)),
	1998 => std_logic_vector(to_unsigned(42, 8)),
	1999 => std_logic_vector(to_unsigned(42, 8)),
	2000 => std_logic_vector(to_unsigned(42, 8)),
	2001 => std_logic_vector(to_unsigned(42, 8)),
	2002 => std_logic_vector(to_unsigned(42, 8)),
	2003 => std_logic_vector(to_unsigned(42, 8)),
	2004 => std_logic_vector(to_unsigned(41, 8)),
	2005 => std_logic_vector(to_unsigned(41, 8)),
	2006 => std_logic_vector(to_unsigned(41, 8)),
	2007 => std_logic_vector(to_unsigned(42, 8)),
	2008 => std_logic_vector(to_unsigned(42, 8)),
	2009 => std_logic_vector(to_unsigned(42, 8)),
	2010 => std_logic_vector(to_unsigned(42, 8)),
	2011 => std_logic_vector(to_unsigned(41, 8)),
	2012 => std_logic_vector(to_unsigned(41, 8)),
	2013 => std_logic_vector(to_unsigned(41, 8)),
	2014 => std_logic_vector(to_unsigned(41, 8)),
	2015 => std_logic_vector(to_unsigned(42, 8)),
	2016 => std_logic_vector(to_unsigned(42, 8)),
	2017 => std_logic_vector(to_unsigned(41, 8)),
	2018 => std_logic_vector(to_unsigned(42, 8)),
	2019 => std_logic_vector(to_unsigned(41, 8)),
	2020 => std_logic_vector(to_unsigned(41, 8)),
	2021 => std_logic_vector(to_unsigned(42, 8)),
	2022 => std_logic_vector(to_unsigned(41, 8)),
	2023 => std_logic_vector(to_unsigned(42, 8)),
	2024 => std_logic_vector(to_unsigned(41, 8)),
	2025 => std_logic_vector(to_unsigned(42, 8)),
	2026 => std_logic_vector(to_unsigned(41, 8)),
	2027 => std_logic_vector(to_unsigned(41, 8)),
	2028 => std_logic_vector(to_unsigned(41, 8)),
	2029 => std_logic_vector(to_unsigned(42, 8)),
	2030 => std_logic_vector(to_unsigned(41, 8)),
	2031 => std_logic_vector(to_unsigned(41, 8)),
	2032 => std_logic_vector(to_unsigned(41, 8)),
	2033 => std_logic_vector(to_unsigned(42, 8)),
	2034 => std_logic_vector(to_unsigned(42, 8)),
	2035 => std_logic_vector(to_unsigned(42, 8)),
	2036 => std_logic_vector(to_unsigned(41, 8)),
	2037 => std_logic_vector(to_unsigned(42, 8)),
	2038 => std_logic_vector(to_unsigned(41, 8)),
	2039 => std_logic_vector(to_unsigned(42, 8)),
	2040 => std_logic_vector(to_unsigned(42, 8)),
	2041 => std_logic_vector(to_unsigned(42, 8)),
	2042 => std_logic_vector(to_unsigned(41, 8)),
	2043 => std_logic_vector(to_unsigned(41, 8)),
	2044 => std_logic_vector(to_unsigned(42, 8)),
	2045 => std_logic_vector(to_unsigned(42, 8)),
	2046 => std_logic_vector(to_unsigned(42, 8)),
	2047 => std_logic_vector(to_unsigned(42, 8)),
	2048 => std_logic_vector(to_unsigned(42, 8)),
	2049 => std_logic_vector(to_unsigned(41, 8)),
	2050 => std_logic_vector(to_unsigned(42, 8)),
	2051 => std_logic_vector(to_unsigned(42, 8)),
	2052 => std_logic_vector(to_unsigned(41, 8)),
	2053 => std_logic_vector(to_unsigned(42, 8)),
	2054 => std_logic_vector(to_unsigned(42, 8)),
	2055 => std_logic_vector(to_unsigned(41, 8)),
	2056 => std_logic_vector(to_unsigned(42, 8)),
	2057 => std_logic_vector(to_unsigned(42, 8)),
	2058 => std_logic_vector(to_unsigned(41, 8)),
	2059 => std_logic_vector(to_unsigned(41, 8)),
	2060 => std_logic_vector(to_unsigned(41, 8)),
	2061 => std_logic_vector(to_unsigned(42, 8)),
	2062 => std_logic_vector(to_unsigned(42, 8)),
	2063 => std_logic_vector(to_unsigned(41, 8)),
	2064 => std_logic_vector(to_unsigned(42, 8)),
	2065 => std_logic_vector(to_unsigned(42, 8)),
	2066 => std_logic_vector(to_unsigned(42, 8)),
	2067 => std_logic_vector(to_unsigned(42, 8)),
	2068 => std_logic_vector(to_unsigned(42, 8)),
	2069 => std_logic_vector(to_unsigned(41, 8)),
	2070 => std_logic_vector(to_unsigned(42, 8)),
	2071 => std_logic_vector(to_unsigned(42, 8)),
	2072 => std_logic_vector(to_unsigned(41, 8)),
	2073 => std_logic_vector(to_unsigned(41, 8)),
	2074 => std_logic_vector(to_unsigned(42, 8)),
	2075 => std_logic_vector(to_unsigned(42, 8)),
	2076 => std_logic_vector(to_unsigned(42, 8)),
	2077 => std_logic_vector(to_unsigned(42, 8)),
	2078 => std_logic_vector(to_unsigned(41, 8)),
	2079 => std_logic_vector(to_unsigned(42, 8)),
	2080 => std_logic_vector(to_unsigned(42, 8)),
	2081 => std_logic_vector(to_unsigned(42, 8)),
	2082 => std_logic_vector(to_unsigned(42, 8)),
	2083 => std_logic_vector(to_unsigned(41, 8)),
	2084 => std_logic_vector(to_unsigned(41, 8)),
	2085 => std_logic_vector(to_unsigned(42, 8)),
	2086 => std_logic_vector(to_unsigned(41, 8)),
	2087 => std_logic_vector(to_unsigned(41, 8)),
	2088 => std_logic_vector(to_unsigned(41, 8)),
	2089 => std_logic_vector(to_unsigned(41, 8)),
	2090 => std_logic_vector(to_unsigned(42, 8)),
	2091 => std_logic_vector(to_unsigned(41, 8)),
	2092 => std_logic_vector(to_unsigned(42, 8)),
	2093 => std_logic_vector(to_unsigned(42, 8)),
	2094 => std_logic_vector(to_unsigned(42, 8)),
	2095 => std_logic_vector(to_unsigned(42, 8)),
	2096 => std_logic_vector(to_unsigned(42, 8)),
	2097 => std_logic_vector(to_unsigned(42, 8)),
	2098 => std_logic_vector(to_unsigned(42, 8)),
	2099 => std_logic_vector(to_unsigned(42, 8)),
	2100 => std_logic_vector(to_unsigned(41, 8)),
	2101 => std_logic_vector(to_unsigned(41, 8)),
	2102 => std_logic_vector(to_unsigned(41, 8)),
	2103 => std_logic_vector(to_unsigned(41, 8)),
	2104 => std_logic_vector(to_unsigned(41, 8)),
	2105 => std_logic_vector(to_unsigned(41, 8)),
	2106 => std_logic_vector(to_unsigned(42, 8)),
	2107 => std_logic_vector(to_unsigned(42, 8)),
	2108 => std_logic_vector(to_unsigned(41, 8)),
	2109 => std_logic_vector(to_unsigned(42, 8)),
	2110 => std_logic_vector(to_unsigned(42, 8)),
	2111 => std_logic_vector(to_unsigned(42, 8)),
	2112 => std_logic_vector(to_unsigned(42, 8)),
	2113 => std_logic_vector(to_unsigned(41, 8)),
	2114 => std_logic_vector(to_unsigned(42, 8)),
	2115 => std_logic_vector(to_unsigned(41, 8)),
	2116 => std_logic_vector(to_unsigned(41, 8)),
	2117 => std_logic_vector(to_unsigned(41, 8)),
	2118 => std_logic_vector(to_unsigned(41, 8)),
	2119 => std_logic_vector(to_unsigned(41, 8)),
	2120 => std_logic_vector(to_unsigned(41, 8)),
	2121 => std_logic_vector(to_unsigned(42, 8)),
	2122 => std_logic_vector(to_unsigned(42, 8)),
	2123 => std_logic_vector(to_unsigned(41, 8)),
	2124 => std_logic_vector(to_unsigned(41, 8)),
	2125 => std_logic_vector(to_unsigned(41, 8)),
	2126 => std_logic_vector(to_unsigned(42, 8)),
	2127 => std_logic_vector(to_unsigned(42, 8)),
	2128 => std_logic_vector(to_unsigned(41, 8)),
	2129 => std_logic_vector(to_unsigned(41, 8)),
	2130 => std_logic_vector(to_unsigned(42, 8)),
	2131 => std_logic_vector(to_unsigned(42, 8)),
	2132 => std_logic_vector(to_unsigned(41, 8)),
	2133 => std_logic_vector(to_unsigned(42, 8)),
	2134 => std_logic_vector(to_unsigned(42, 8)),
	2135 => std_logic_vector(to_unsigned(42, 8)),
	2136 => std_logic_vector(to_unsigned(42, 8)),
	2137 => std_logic_vector(to_unsigned(42, 8)),
	2138 => std_logic_vector(to_unsigned(41, 8)),
	2139 => std_logic_vector(to_unsigned(41, 8)),
	2140 => std_logic_vector(to_unsigned(42, 8)),
	2141 => std_logic_vector(to_unsigned(41, 8)),
	2142 => std_logic_vector(to_unsigned(41, 8)),
	2143 => std_logic_vector(to_unsigned(42, 8)),
	2144 => std_logic_vector(to_unsigned(41, 8)),
	2145 => std_logic_vector(to_unsigned(41, 8)),
	2146 => std_logic_vector(to_unsigned(41, 8)),
	2147 => std_logic_vector(to_unsigned(42, 8)),
	2148 => std_logic_vector(to_unsigned(41, 8)),
	2149 => std_logic_vector(to_unsigned(42, 8)),
	2150 => std_logic_vector(to_unsigned(42, 8)),
	2151 => std_logic_vector(to_unsigned(42, 8)),
	2152 => std_logic_vector(to_unsigned(42, 8)),
	2153 => std_logic_vector(to_unsigned(42, 8)),
	2154 => std_logic_vector(to_unsigned(41, 8)),
	2155 => std_logic_vector(to_unsigned(41, 8)),
	2156 => std_logic_vector(to_unsigned(42, 8)),
	2157 => std_logic_vector(to_unsigned(41, 8)),
	2158 => std_logic_vector(to_unsigned(42, 8)),
	2159 => std_logic_vector(to_unsigned(42, 8)),
	2160 => std_logic_vector(to_unsigned(42, 8)),
	2161 => std_logic_vector(to_unsigned(42, 8)),
	2162 => std_logic_vector(to_unsigned(41, 8)),
	2163 => std_logic_vector(to_unsigned(41, 8)),
	2164 => std_logic_vector(to_unsigned(42, 8)),
	2165 => std_logic_vector(to_unsigned(41, 8)),
	2166 => std_logic_vector(to_unsigned(41, 8)),
	2167 => std_logic_vector(to_unsigned(42, 8)),
	2168 => std_logic_vector(to_unsigned(41, 8)),
	2169 => std_logic_vector(to_unsigned(42, 8)),
	2170 => std_logic_vector(to_unsigned(41, 8)),
	2171 => std_logic_vector(to_unsigned(42, 8)),
	2172 => std_logic_vector(to_unsigned(41, 8)),
	2173 => std_logic_vector(to_unsigned(41, 8)),
	2174 => std_logic_vector(to_unsigned(42, 8)),
	2175 => std_logic_vector(to_unsigned(42, 8)),
	2176 => std_logic_vector(to_unsigned(41, 8)),
	2177 => std_logic_vector(to_unsigned(41, 8)),
	2178 => std_logic_vector(to_unsigned(41, 8)),
	2179 => std_logic_vector(to_unsigned(42, 8)),
	2180 => std_logic_vector(to_unsigned(41, 8)),
	2181 => std_logic_vector(to_unsigned(42, 8)),
	2182 => std_logic_vector(to_unsigned(41, 8)),
	2183 => std_logic_vector(to_unsigned(41, 8)),
	2184 => std_logic_vector(to_unsigned(42, 8)),
	2185 => std_logic_vector(to_unsigned(41, 8)),
	2186 => std_logic_vector(to_unsigned(41, 8)),
	2187 => std_logic_vector(to_unsigned(42, 8)),
	2188 => std_logic_vector(to_unsigned(41, 8)),
	2189 => std_logic_vector(to_unsigned(41, 8)),
	2190 => std_logic_vector(to_unsigned(42, 8)),
	2191 => std_logic_vector(to_unsigned(41, 8)),
	2192 => std_logic_vector(to_unsigned(42, 8)),
	2193 => std_logic_vector(to_unsigned(42, 8)),
	2194 => std_logic_vector(to_unsigned(41, 8)),
	2195 => std_logic_vector(to_unsigned(41, 8)),
	2196 => std_logic_vector(to_unsigned(42, 8)),
	2197 => std_logic_vector(to_unsigned(41, 8)),
	2198 => std_logic_vector(to_unsigned(41, 8)),
	2199 => std_logic_vector(to_unsigned(42, 8)),
	2200 => std_logic_vector(to_unsigned(41, 8)),
	2201 => std_logic_vector(to_unsigned(41, 8)),
	2202 => std_logic_vector(to_unsigned(42, 8)),
	2203 => std_logic_vector(to_unsigned(42, 8)),
	2204 => std_logic_vector(to_unsigned(41, 8)),
	2205 => std_logic_vector(to_unsigned(42, 8)),
	2206 => std_logic_vector(to_unsigned(41, 8)),
	2207 => std_logic_vector(to_unsigned(42, 8)),
	2208 => std_logic_vector(to_unsigned(42, 8)),
	2209 => std_logic_vector(to_unsigned(42, 8)),
	2210 => std_logic_vector(to_unsigned(42, 8)),
	2211 => std_logic_vector(to_unsigned(41, 8)),
	2212 => std_logic_vector(to_unsigned(41, 8)),
	2213 => std_logic_vector(to_unsigned(42, 8)),
	2214 => std_logic_vector(to_unsigned(42, 8)),
	2215 => std_logic_vector(to_unsigned(42, 8)),
	2216 => std_logic_vector(to_unsigned(42, 8)),
	2217 => std_logic_vector(to_unsigned(42, 8)),
	2218 => std_logic_vector(to_unsigned(41, 8)),
	2219 => std_logic_vector(to_unsigned(41, 8)),
	2220 => std_logic_vector(to_unsigned(41, 8)),
	2221 => std_logic_vector(to_unsigned(41, 8)),
	2222 => std_logic_vector(to_unsigned(41, 8)),
	2223 => std_logic_vector(to_unsigned(41, 8)),
	2224 => std_logic_vector(to_unsigned(42, 8)),
	2225 => std_logic_vector(to_unsigned(42, 8)),
	2226 => std_logic_vector(to_unsigned(42, 8)),
	2227 => std_logic_vector(to_unsigned(41, 8)),
	2228 => std_logic_vector(to_unsigned(42, 8)),
	2229 => std_logic_vector(to_unsigned(41, 8)),
	2230 => std_logic_vector(to_unsigned(41, 8)),
	2231 => std_logic_vector(to_unsigned(41, 8)),
	2232 => std_logic_vector(to_unsigned(42, 8)),
	2233 => std_logic_vector(to_unsigned(42, 8)),
	2234 => std_logic_vector(to_unsigned(41, 8)),
	2235 => std_logic_vector(to_unsigned(41, 8)),
	2236 => std_logic_vector(to_unsigned(42, 8)),
	2237 => std_logic_vector(to_unsigned(42, 8)),
	2238 => std_logic_vector(to_unsigned(41, 8)),
	2239 => std_logic_vector(to_unsigned(42, 8)),
	2240 => std_logic_vector(to_unsigned(42, 8)),
	2241 => std_logic_vector(to_unsigned(41, 8)),
	2242 => std_logic_vector(to_unsigned(41, 8)),
	2243 => std_logic_vector(to_unsigned(41, 8)),
	2244 => std_logic_vector(to_unsigned(42, 8)),
	2245 => std_logic_vector(to_unsigned(41, 8)),
	2246 => std_logic_vector(to_unsigned(42, 8)),
	2247 => std_logic_vector(to_unsigned(41, 8)),
	2248 => std_logic_vector(to_unsigned(42, 8)),
	2249 => std_logic_vector(to_unsigned(42, 8)),
	2250 => std_logic_vector(to_unsigned(42, 8)),
	2251 => std_logic_vector(to_unsigned(41, 8)),
	2252 => std_logic_vector(to_unsigned(41, 8)),
	2253 => std_logic_vector(to_unsigned(41, 8)),
	2254 => std_logic_vector(to_unsigned(42, 8)),
	2255 => std_logic_vector(to_unsigned(42, 8)),
	2256 => std_logic_vector(to_unsigned(42, 8)),
	2257 => std_logic_vector(to_unsigned(42, 8)),
	2258 => std_logic_vector(to_unsigned(42, 8)),
	2259 => std_logic_vector(to_unsigned(41, 8)),
	2260 => std_logic_vector(to_unsigned(41, 8)),
	2261 => std_logic_vector(to_unsigned(41, 8)),
	2262 => std_logic_vector(to_unsigned(41, 8)),
	2263 => std_logic_vector(to_unsigned(42, 8)),
	2264 => std_logic_vector(to_unsigned(41, 8)),
	2265 => std_logic_vector(to_unsigned(42, 8)),
	2266 => std_logic_vector(to_unsigned(41, 8)),
	2267 => std_logic_vector(to_unsigned(41, 8)),
	2268 => std_logic_vector(to_unsigned(41, 8)),
	2269 => std_logic_vector(to_unsigned(41, 8)),
	2270 => std_logic_vector(to_unsigned(41, 8)),
	2271 => std_logic_vector(to_unsigned(41, 8)),
	2272 => std_logic_vector(to_unsigned(42, 8)),
	2273 => std_logic_vector(to_unsigned(41, 8)),
	2274 => std_logic_vector(to_unsigned(41, 8)),
	2275 => std_logic_vector(to_unsigned(41, 8)),
	2276 => std_logic_vector(to_unsigned(42, 8)),
	2277 => std_logic_vector(to_unsigned(41, 8)),
	2278 => std_logic_vector(to_unsigned(42, 8)),
	2279 => std_logic_vector(to_unsigned(41, 8)),
	2280 => std_logic_vector(to_unsigned(42, 8)),
	2281 => std_logic_vector(to_unsigned(42, 8)),
	2282 => std_logic_vector(to_unsigned(41, 8)),
	2283 => std_logic_vector(to_unsigned(42, 8)),
	2284 => std_logic_vector(to_unsigned(42, 8)),
	2285 => std_logic_vector(to_unsigned(41, 8)),
	2286 => std_logic_vector(to_unsigned(41, 8)),
	2287 => std_logic_vector(to_unsigned(42, 8)),
	2288 => std_logic_vector(to_unsigned(41, 8)),
	2289 => std_logic_vector(to_unsigned(41, 8)),
	2290 => std_logic_vector(to_unsigned(41, 8)),
	2291 => std_logic_vector(to_unsigned(42, 8)),
	2292 => std_logic_vector(to_unsigned(42, 8)),
	2293 => std_logic_vector(to_unsigned(41, 8)),
	2294 => std_logic_vector(to_unsigned(42, 8)),
	2295 => std_logic_vector(to_unsigned(41, 8)),
	2296 => std_logic_vector(to_unsigned(42, 8)),
	2297 => std_logic_vector(to_unsigned(42, 8)),
	2298 => std_logic_vector(to_unsigned(41, 8)),
	2299 => std_logic_vector(to_unsigned(42, 8)),
	2300 => std_logic_vector(to_unsigned(42, 8)),
	2301 => std_logic_vector(to_unsigned(41, 8)),
	2302 => std_logic_vector(to_unsigned(42, 8)),
	2303 => std_logic_vector(to_unsigned(41, 8)),
	2304 => std_logic_vector(to_unsigned(42, 8)),
	2305 => std_logic_vector(to_unsigned(41, 8)),
	2306 => std_logic_vector(to_unsigned(42, 8)),
	2307 => std_logic_vector(to_unsigned(41, 8)),
	2308 => std_logic_vector(to_unsigned(42, 8)),
	2309 => std_logic_vector(to_unsigned(42, 8)),
	2310 => std_logic_vector(to_unsigned(42, 8)),
	2311 => std_logic_vector(to_unsigned(42, 8)),
	2312 => std_logic_vector(to_unsigned(42, 8)),
	2313 => std_logic_vector(to_unsigned(42, 8)),
	2314 => std_logic_vector(to_unsigned(41, 8)),
	2315 => std_logic_vector(to_unsigned(42, 8)),
	2316 => std_logic_vector(to_unsigned(41, 8)),
	2317 => std_logic_vector(to_unsigned(41, 8)),
	2318 => std_logic_vector(to_unsigned(42, 8)),
	2319 => std_logic_vector(to_unsigned(41, 8)),
	2320 => std_logic_vector(to_unsigned(41, 8)),
	2321 => std_logic_vector(to_unsigned(42, 8)),
	2322 => std_logic_vector(to_unsigned(41, 8)),
	2323 => std_logic_vector(to_unsigned(42, 8)),
	2324 => std_logic_vector(to_unsigned(42, 8)),
	2325 => std_logic_vector(to_unsigned(42, 8)),
	2326 => std_logic_vector(to_unsigned(41, 8)),
	2327 => std_logic_vector(to_unsigned(41, 8)),
	2328 => std_logic_vector(to_unsigned(42, 8)),
	2329 => std_logic_vector(to_unsigned(42, 8)),
	2330 => std_logic_vector(to_unsigned(42, 8)),
	2331 => std_logic_vector(to_unsigned(42, 8)),
	2332 => std_logic_vector(to_unsigned(41, 8)),
	2333 => std_logic_vector(to_unsigned(42, 8)),
	2334 => std_logic_vector(to_unsigned(42, 8)),
	2335 => std_logic_vector(to_unsigned(42, 8)),
	2336 => std_logic_vector(to_unsigned(41, 8)),
	2337 => std_logic_vector(to_unsigned(41, 8)),
	2338 => std_logic_vector(to_unsigned(42, 8)),
	2339 => std_logic_vector(to_unsigned(42, 8)),
	2340 => std_logic_vector(to_unsigned(41, 8)),
	2341 => std_logic_vector(to_unsigned(42, 8)),
	2342 => std_logic_vector(to_unsigned(41, 8)),
	2343 => std_logic_vector(to_unsigned(41, 8)),
	2344 => std_logic_vector(to_unsigned(41, 8)),
	2345 => std_logic_vector(to_unsigned(42, 8)),
	2346 => std_logic_vector(to_unsigned(42, 8)),
	2347 => std_logic_vector(to_unsigned(41, 8)),
	2348 => std_logic_vector(to_unsigned(42, 8)),
	2349 => std_logic_vector(to_unsigned(41, 8)),
	2350 => std_logic_vector(to_unsigned(42, 8)),
	2351 => std_logic_vector(to_unsigned(41, 8)),
	2352 => std_logic_vector(to_unsigned(42, 8)),
	2353 => std_logic_vector(to_unsigned(41, 8)),
	2354 => std_logic_vector(to_unsigned(41, 8)),
	2355 => std_logic_vector(to_unsigned(41, 8)),
	2356 => std_logic_vector(to_unsigned(41, 8)),
	2357 => std_logic_vector(to_unsigned(41, 8)),
	2358 => std_logic_vector(to_unsigned(41, 8)),
	2359 => std_logic_vector(to_unsigned(42, 8)),
	2360 => std_logic_vector(to_unsigned(41, 8)),
	2361 => std_logic_vector(to_unsigned(41, 8)),
	2362 => std_logic_vector(to_unsigned(42, 8)),
	2363 => std_logic_vector(to_unsigned(42, 8)),
	2364 => std_logic_vector(to_unsigned(42, 8)),
	2365 => std_logic_vector(to_unsigned(41, 8)),
	2366 => std_logic_vector(to_unsigned(41, 8)),
	2367 => std_logic_vector(to_unsigned(41, 8)),
	2368 => std_logic_vector(to_unsigned(42, 8)),
	2369 => std_logic_vector(to_unsigned(41, 8)),
	2370 => std_logic_vector(to_unsigned(41, 8)),
	2371 => std_logic_vector(to_unsigned(41, 8)),
	2372 => std_logic_vector(to_unsigned(41, 8)),
	2373 => std_logic_vector(to_unsigned(41, 8)),
	2374 => std_logic_vector(to_unsigned(42, 8)),
	2375 => std_logic_vector(to_unsigned(42, 8)),
	2376 => std_logic_vector(to_unsigned(42, 8)),
	2377 => std_logic_vector(to_unsigned(42, 8)),
	2378 => std_logic_vector(to_unsigned(42, 8)),
	2379 => std_logic_vector(to_unsigned(42, 8)),
	2380 => std_logic_vector(to_unsigned(41, 8)),
	2381 => std_logic_vector(to_unsigned(42, 8)),
	2382 => std_logic_vector(to_unsigned(41, 8)),
	2383 => std_logic_vector(to_unsigned(42, 8)),
	2384 => std_logic_vector(to_unsigned(42, 8)),
	2385 => std_logic_vector(to_unsigned(41, 8)),
	2386 => std_logic_vector(to_unsigned(42, 8)),
	2387 => std_logic_vector(to_unsigned(42, 8)),
	2388 => std_logic_vector(to_unsigned(41, 8)),
	2389 => std_logic_vector(to_unsigned(42, 8)),
	2390 => std_logic_vector(to_unsigned(42, 8)),
	2391 => std_logic_vector(to_unsigned(41, 8)),
	2392 => std_logic_vector(to_unsigned(41, 8)),
	2393 => std_logic_vector(to_unsigned(41, 8)),
	2394 => std_logic_vector(to_unsigned(42, 8)),
	2395 => std_logic_vector(to_unsigned(42, 8)),
	2396 => std_logic_vector(to_unsigned(41, 8)),
	2397 => std_logic_vector(to_unsigned(42, 8)),
	2398 => std_logic_vector(to_unsigned(42, 8)),
	2399 => std_logic_vector(to_unsigned(42, 8)),
	2400 => std_logic_vector(to_unsigned(42, 8)),
	2401 => std_logic_vector(to_unsigned(41, 8)),
	2402 => std_logic_vector(to_unsigned(41, 8)),
	2403 => std_logic_vector(to_unsigned(41, 8)),
	2404 => std_logic_vector(to_unsigned(42, 8)),
	2405 => std_logic_vector(to_unsigned(42, 8)),
	2406 => std_logic_vector(to_unsigned(41, 8)),
	2407 => std_logic_vector(to_unsigned(41, 8)),
	2408 => std_logic_vector(to_unsigned(41, 8)),
	2409 => std_logic_vector(to_unsigned(41, 8)),
	2410 => std_logic_vector(to_unsigned(41, 8)),
	2411 => std_logic_vector(to_unsigned(41, 8)),
	2412 => std_logic_vector(to_unsigned(42, 8)),
	2413 => std_logic_vector(to_unsigned(41, 8)),
	2414 => std_logic_vector(to_unsigned(41, 8)),
	2415 => std_logic_vector(to_unsigned(41, 8)),
	2416 => std_logic_vector(to_unsigned(41, 8)),
	2417 => std_logic_vector(to_unsigned(42, 8)),
	2418 => std_logic_vector(to_unsigned(42, 8)),
	2419 => std_logic_vector(to_unsigned(42, 8)),
	2420 => std_logic_vector(to_unsigned(42, 8)),
	2421 => std_logic_vector(to_unsigned(42, 8)),
	2422 => std_logic_vector(to_unsigned(41, 8)),
	2423 => std_logic_vector(to_unsigned(42, 8)),
	2424 => std_logic_vector(to_unsigned(41, 8)),
	2425 => std_logic_vector(to_unsigned(41, 8)),
	2426 => std_logic_vector(to_unsigned(41, 8)),
	2427 => std_logic_vector(to_unsigned(42, 8)),
	2428 => std_logic_vector(to_unsigned(41, 8)),
	2429 => std_logic_vector(to_unsigned(41, 8)),
	2430 => std_logic_vector(to_unsigned(42, 8)),
	2431 => std_logic_vector(to_unsigned(42, 8)),
	2432 => std_logic_vector(to_unsigned(42, 8)),
	2433 => std_logic_vector(to_unsigned(42, 8)),
	2434 => std_logic_vector(to_unsigned(42, 8)),
	2435 => std_logic_vector(to_unsigned(42, 8)),
	2436 => std_logic_vector(to_unsigned(42, 8)),
	2437 => std_logic_vector(to_unsigned(41, 8)),
	2438 => std_logic_vector(to_unsigned(41, 8)),
	2439 => std_logic_vector(to_unsigned(41, 8)),
	2440 => std_logic_vector(to_unsigned(41, 8)),
	2441 => std_logic_vector(to_unsigned(41, 8)),
	2442 => std_logic_vector(to_unsigned(41, 8)),
	2443 => std_logic_vector(to_unsigned(42, 8)),
	2444 => std_logic_vector(to_unsigned(42, 8)),
	2445 => std_logic_vector(to_unsigned(42, 8)),
	2446 => std_logic_vector(to_unsigned(42, 8)),
	2447 => std_logic_vector(to_unsigned(42, 8)),
	2448 => std_logic_vector(to_unsigned(41, 8)),
	2449 => std_logic_vector(to_unsigned(41, 8)),
	2450 => std_logic_vector(to_unsigned(42, 8)),
	2451 => std_logic_vector(to_unsigned(42, 8)),
	2452 => std_logic_vector(to_unsigned(42, 8)),
	2453 => std_logic_vector(to_unsigned(41, 8)),
	2454 => std_logic_vector(to_unsigned(41, 8)),
	2455 => std_logic_vector(to_unsigned(42, 8)),
	2456 => std_logic_vector(to_unsigned(41, 8)),
	2457 => std_logic_vector(to_unsigned(42, 8)),
	2458 => std_logic_vector(to_unsigned(41, 8)),
	2459 => std_logic_vector(to_unsigned(41, 8)),
	2460 => std_logic_vector(to_unsigned(41, 8)),
	2461 => std_logic_vector(to_unsigned(42, 8)),
	2462 => std_logic_vector(to_unsigned(41, 8)),
	2463 => std_logic_vector(to_unsigned(42, 8)),
	2464 => std_logic_vector(to_unsigned(42, 8)),
	2465 => std_logic_vector(to_unsigned(41, 8)),
	2466 => std_logic_vector(to_unsigned(41, 8)),
	2467 => std_logic_vector(to_unsigned(42, 8)),
	2468 => std_logic_vector(to_unsigned(42, 8)),
	2469 => std_logic_vector(to_unsigned(41, 8)),
	2470 => std_logic_vector(to_unsigned(42, 8)),
	2471 => std_logic_vector(to_unsigned(41, 8)),
	2472 => std_logic_vector(to_unsigned(41, 8)),
	2473 => std_logic_vector(to_unsigned(41, 8)),
	2474 => std_logic_vector(to_unsigned(41, 8)),
	2475 => std_logic_vector(to_unsigned(42, 8)),
	2476 => std_logic_vector(to_unsigned(42, 8)),
	2477 => std_logic_vector(to_unsigned(42, 8)),
	2478 => std_logic_vector(to_unsigned(42, 8)),
	2479 => std_logic_vector(to_unsigned(42, 8)),
	2480 => std_logic_vector(to_unsigned(42, 8)),
	2481 => std_logic_vector(to_unsigned(42, 8)),
	2482 => std_logic_vector(to_unsigned(41, 8)),
	2483 => std_logic_vector(to_unsigned(41, 8)),
	2484 => std_logic_vector(to_unsigned(41, 8)),
	2485 => std_logic_vector(to_unsigned(41, 8)),
	2486 => std_logic_vector(to_unsigned(41, 8)),
	2487 => std_logic_vector(to_unsigned(42, 8)),
	2488 => std_logic_vector(to_unsigned(41, 8)),
	2489 => std_logic_vector(to_unsigned(41, 8)),
	2490 => std_logic_vector(to_unsigned(42, 8)),
	2491 => std_logic_vector(to_unsigned(42, 8)),
	2492 => std_logic_vector(to_unsigned(42, 8)),
	2493 => std_logic_vector(to_unsigned(42, 8)),
	2494 => std_logic_vector(to_unsigned(41, 8)),
	2495 => std_logic_vector(to_unsigned(41, 8)),
	2496 => std_logic_vector(to_unsigned(42, 8)),
	2497 => std_logic_vector(to_unsigned(41, 8)),
	2498 => std_logic_vector(to_unsigned(42, 8)),
	2499 => std_logic_vector(to_unsigned(41, 8)),
	2500 => std_logic_vector(to_unsigned(42, 8)),
	2501 => std_logic_vector(to_unsigned(41, 8)),
	2502 => std_logic_vector(to_unsigned(42, 8)),
	2503 => std_logic_vector(to_unsigned(41, 8)),
	2504 => std_logic_vector(to_unsigned(42, 8)),
	2505 => std_logic_vector(to_unsigned(41, 8)),
	2506 => std_logic_vector(to_unsigned(41, 8)),
	2507 => std_logic_vector(to_unsigned(42, 8)),
	2508 => std_logic_vector(to_unsigned(42, 8)),
	2509 => std_logic_vector(to_unsigned(42, 8)),
	2510 => std_logic_vector(to_unsigned(41, 8)),
	2511 => std_logic_vector(to_unsigned(41, 8)),
	2512 => std_logic_vector(to_unsigned(42, 8)),
	2513 => std_logic_vector(to_unsigned(41, 8)),
	2514 => std_logic_vector(to_unsigned(41, 8)),
	2515 => std_logic_vector(to_unsigned(42, 8)),
	2516 => std_logic_vector(to_unsigned(42, 8)),
	2517 => std_logic_vector(to_unsigned(42, 8)),
	2518 => std_logic_vector(to_unsigned(41, 8)),
	2519 => std_logic_vector(to_unsigned(42, 8)),
	2520 => std_logic_vector(to_unsigned(42, 8)),
	2521 => std_logic_vector(to_unsigned(41, 8)),
	2522 => std_logic_vector(to_unsigned(41, 8)),
	2523 => std_logic_vector(to_unsigned(41, 8)),
	2524 => std_logic_vector(to_unsigned(42, 8)),
	2525 => std_logic_vector(to_unsigned(42, 8)),
	2526 => std_logic_vector(to_unsigned(41, 8)),
	2527 => std_logic_vector(to_unsigned(41, 8)),
	2528 => std_logic_vector(to_unsigned(42, 8)),
	2529 => std_logic_vector(to_unsigned(41, 8)),
	2530 => std_logic_vector(to_unsigned(42, 8)),
	2531 => std_logic_vector(to_unsigned(42, 8)),
	2532 => std_logic_vector(to_unsigned(42, 8)),
	2533 => std_logic_vector(to_unsigned(41, 8)),
	2534 => std_logic_vector(to_unsigned(41, 8)),
	2535 => std_logic_vector(to_unsigned(41, 8)),
	2536 => std_logic_vector(to_unsigned(42, 8)),
	2537 => std_logic_vector(to_unsigned(42, 8)),
	2538 => std_logic_vector(to_unsigned(41, 8)),
	2539 => std_logic_vector(to_unsigned(42, 8)),
	2540 => std_logic_vector(to_unsigned(41, 8)),
	2541 => std_logic_vector(to_unsigned(41, 8)),
	2542 => std_logic_vector(to_unsigned(42, 8)),
	2543 => std_logic_vector(to_unsigned(41, 8)),
	2544 => std_logic_vector(to_unsigned(42, 8)),
	2545 => std_logic_vector(to_unsigned(42, 8)),
	2546 => std_logic_vector(to_unsigned(41, 8)),
	2547 => std_logic_vector(to_unsigned(42, 8)),
	2548 => std_logic_vector(to_unsigned(41, 8)),
	2549 => std_logic_vector(to_unsigned(41, 8)),
	2550 => std_logic_vector(to_unsigned(42, 8)),
	2551 => std_logic_vector(to_unsigned(42, 8)),
	2552 => std_logic_vector(to_unsigned(42, 8)),
	2553 => std_logic_vector(to_unsigned(41, 8)),
	2554 => std_logic_vector(to_unsigned(42, 8)),
	2555 => std_logic_vector(to_unsigned(42, 8)),
	2556 => std_logic_vector(to_unsigned(41, 8)),
	2557 => std_logic_vector(to_unsigned(42, 8)),
	2558 => std_logic_vector(to_unsigned(42, 8)),
	2559 => std_logic_vector(to_unsigned(42, 8)),
	2560 => std_logic_vector(to_unsigned(41, 8)),
	2561 => std_logic_vector(to_unsigned(41, 8)),
	2562 => std_logic_vector(to_unsigned(42, 8)),
	2563 => std_logic_vector(to_unsigned(41, 8)),
	2564 => std_logic_vector(to_unsigned(42, 8)),
	2565 => std_logic_vector(to_unsigned(42, 8)),
	2566 => std_logic_vector(to_unsigned(42, 8)),
	2567 => std_logic_vector(to_unsigned(42, 8)),
	2568 => std_logic_vector(to_unsigned(42, 8)),
	2569 => std_logic_vector(to_unsigned(41, 8)),
	2570 => std_logic_vector(to_unsigned(41, 8)),
	2571 => std_logic_vector(to_unsigned(42, 8)),
	2572 => std_logic_vector(to_unsigned(42, 8)),
	2573 => std_logic_vector(to_unsigned(41, 8)),
	2574 => std_logic_vector(to_unsigned(41, 8)),
	2575 => std_logic_vector(to_unsigned(41, 8)),
	2576 => std_logic_vector(to_unsigned(41, 8)),
	2577 => std_logic_vector(to_unsigned(42, 8)),
	2578 => std_logic_vector(to_unsigned(42, 8)),
	2579 => std_logic_vector(to_unsigned(41, 8)),
	2580 => std_logic_vector(to_unsigned(41, 8)),
	2581 => std_logic_vector(to_unsigned(41, 8)),
	2582 => std_logic_vector(to_unsigned(41, 8)),
	2583 => std_logic_vector(to_unsigned(42, 8)),
	2584 => std_logic_vector(to_unsigned(42, 8)),
	2585 => std_logic_vector(to_unsigned(42, 8)),
	2586 => std_logic_vector(to_unsigned(41, 8)),
	2587 => std_logic_vector(to_unsigned(42, 8)),
	2588 => std_logic_vector(to_unsigned(42, 8)),
	2589 => std_logic_vector(to_unsigned(42, 8)),
	2590 => std_logic_vector(to_unsigned(42, 8)),
	2591 => std_logic_vector(to_unsigned(41, 8)),
	2592 => std_logic_vector(to_unsigned(41, 8)),
	2593 => std_logic_vector(to_unsigned(42, 8)),
	2594 => std_logic_vector(to_unsigned(42, 8)),
	2595 => std_logic_vector(to_unsigned(41, 8)),
	2596 => std_logic_vector(to_unsigned(41, 8)),
	2597 => std_logic_vector(to_unsigned(41, 8)),
	2598 => std_logic_vector(to_unsigned(42, 8)),
	2599 => std_logic_vector(to_unsigned(42, 8)),
	2600 => std_logic_vector(to_unsigned(41, 8)),
	2601 => std_logic_vector(to_unsigned(41, 8)),
	2602 => std_logic_vector(to_unsigned(42, 8)),
	2603 => std_logic_vector(to_unsigned(42, 8)),
	2604 => std_logic_vector(to_unsigned(42, 8)),
	2605 => std_logic_vector(to_unsigned(42, 8)),
	2606 => std_logic_vector(to_unsigned(42, 8)),
	2607 => std_logic_vector(to_unsigned(41, 8)),
	2608 => std_logic_vector(to_unsigned(41, 8)),
	2609 => std_logic_vector(to_unsigned(41, 8)),
	2610 => std_logic_vector(to_unsigned(42, 8)),
	2611 => std_logic_vector(to_unsigned(42, 8)),
	2612 => std_logic_vector(to_unsigned(41, 8)),
	2613 => std_logic_vector(to_unsigned(41, 8)),
	2614 => std_logic_vector(to_unsigned(42, 8)),
	2615 => std_logic_vector(to_unsigned(42, 8)),
	2616 => std_logic_vector(to_unsigned(41, 8)),
	2617 => std_logic_vector(to_unsigned(41, 8)),
	2618 => std_logic_vector(to_unsigned(41, 8)),
	2619 => std_logic_vector(to_unsigned(42, 8)),
	2620 => std_logic_vector(to_unsigned(41, 8)),
	2621 => std_logic_vector(to_unsigned(42, 8)),
	2622 => std_logic_vector(to_unsigned(42, 8)),
	2623 => std_logic_vector(to_unsigned(42, 8)),
	2624 => std_logic_vector(to_unsigned(41, 8)),
	2625 => std_logic_vector(to_unsigned(42, 8)),
	2626 => std_logic_vector(to_unsigned(42, 8)),
	2627 => std_logic_vector(to_unsigned(41, 8)),
	2628 => std_logic_vector(to_unsigned(42, 8)),
	2629 => std_logic_vector(to_unsigned(41, 8)),
	2630 => std_logic_vector(to_unsigned(41, 8)),
	2631 => std_logic_vector(to_unsigned(41, 8)),
	2632 => std_logic_vector(to_unsigned(42, 8)),
	2633 => std_logic_vector(to_unsigned(41, 8)),
	2634 => std_logic_vector(to_unsigned(41, 8)),
	2635 => std_logic_vector(to_unsigned(41, 8)),
	2636 => std_logic_vector(to_unsigned(42, 8)),
	2637 => std_logic_vector(to_unsigned(42, 8)),
	2638 => std_logic_vector(to_unsigned(42, 8)),
	2639 => std_logic_vector(to_unsigned(42, 8)),
	2640 => std_logic_vector(to_unsigned(42, 8)),
	2641 => std_logic_vector(to_unsigned(41, 8)),
	2642 => std_logic_vector(to_unsigned(42, 8)),
	2643 => std_logic_vector(to_unsigned(41, 8)),
	2644 => std_logic_vector(to_unsigned(42, 8)),
	2645 => std_logic_vector(to_unsigned(42, 8)),
	2646 => std_logic_vector(to_unsigned(41, 8)),
	2647 => std_logic_vector(to_unsigned(42, 8)),
	2648 => std_logic_vector(to_unsigned(41, 8)),
	2649 => std_logic_vector(to_unsigned(42, 8)),
	2650 => std_logic_vector(to_unsigned(42, 8)),
	2651 => std_logic_vector(to_unsigned(42, 8)),
	2652 => std_logic_vector(to_unsigned(41, 8)),
	2653 => std_logic_vector(to_unsigned(41, 8)),
	2654 => std_logic_vector(to_unsigned(41, 8)),
	2655 => std_logic_vector(to_unsigned(42, 8)),
	2656 => std_logic_vector(to_unsigned(41, 8)),
	2657 => std_logic_vector(to_unsigned(41, 8)),
	2658 => std_logic_vector(to_unsigned(41, 8)),
	2659 => std_logic_vector(to_unsigned(42, 8)),
	2660 => std_logic_vector(to_unsigned(42, 8)),
	2661 => std_logic_vector(to_unsigned(42, 8)),
	2662 => std_logic_vector(to_unsigned(41, 8)),
	2663 => std_logic_vector(to_unsigned(41, 8)),
	2664 => std_logic_vector(to_unsigned(42, 8)),
	2665 => std_logic_vector(to_unsigned(41, 8)),
	2666 => std_logic_vector(to_unsigned(41, 8)),
	2667 => std_logic_vector(to_unsigned(42, 8)),
	2668 => std_logic_vector(to_unsigned(42, 8)),
	2669 => std_logic_vector(to_unsigned(41, 8)),
	2670 => std_logic_vector(to_unsigned(42, 8)),
	2671 => std_logic_vector(to_unsigned(42, 8)),
	2672 => std_logic_vector(to_unsigned(41, 8)),
	2673 => std_logic_vector(to_unsigned(42, 8)),
	2674 => std_logic_vector(to_unsigned(41, 8)),
	2675 => std_logic_vector(to_unsigned(42, 8)),
	2676 => std_logic_vector(to_unsigned(41, 8)),
	2677 => std_logic_vector(to_unsigned(41, 8)),
	2678 => std_logic_vector(to_unsigned(42, 8)),
	2679 => std_logic_vector(to_unsigned(41, 8)),
	2680 => std_logic_vector(to_unsigned(42, 8)),
	2681 => std_logic_vector(to_unsigned(41, 8)),
	2682 => std_logic_vector(to_unsigned(41, 8)),
	2683 => std_logic_vector(to_unsigned(42, 8)),
	2684 => std_logic_vector(to_unsigned(41, 8)),
	2685 => std_logic_vector(to_unsigned(41, 8)),
	2686 => std_logic_vector(to_unsigned(42, 8)),
	2687 => std_logic_vector(to_unsigned(41, 8)),
	2688 => std_logic_vector(to_unsigned(41, 8)),
	2689 => std_logic_vector(to_unsigned(42, 8)),
	2690 => std_logic_vector(to_unsigned(42, 8)),
	2691 => std_logic_vector(to_unsigned(42, 8)),
	2692 => std_logic_vector(to_unsigned(42, 8)),
	2693 => std_logic_vector(to_unsigned(42, 8)),
	2694 => std_logic_vector(to_unsigned(41, 8)),
	2695 => std_logic_vector(to_unsigned(42, 8)),
	2696 => std_logic_vector(to_unsigned(41, 8)),
	2697 => std_logic_vector(to_unsigned(42, 8)),
	2698 => std_logic_vector(to_unsigned(41, 8)),
	2699 => std_logic_vector(to_unsigned(42, 8)),
	2700 => std_logic_vector(to_unsigned(41, 8)),
	2701 => std_logic_vector(to_unsigned(42, 8)),
	2702 => std_logic_vector(to_unsigned(42, 8)),
	2703 => std_logic_vector(to_unsigned(41, 8)),
	2704 => std_logic_vector(to_unsigned(42, 8)),
	2705 => std_logic_vector(to_unsigned(42, 8)),
	2706 => std_logic_vector(to_unsigned(42, 8)),
	2707 => std_logic_vector(to_unsigned(42, 8)),
	2708 => std_logic_vector(to_unsigned(42, 8)),
	2709 => std_logic_vector(to_unsigned(41, 8)),
	2710 => std_logic_vector(to_unsigned(41, 8)),
	2711 => std_logic_vector(to_unsigned(42, 8)),
	2712 => std_logic_vector(to_unsigned(41, 8)),
	2713 => std_logic_vector(to_unsigned(41, 8)),
	2714 => std_logic_vector(to_unsigned(41, 8)),
	2715 => std_logic_vector(to_unsigned(42, 8)),
	2716 => std_logic_vector(to_unsigned(42, 8)),
	2717 => std_logic_vector(to_unsigned(41, 8)),
	2718 => std_logic_vector(to_unsigned(41, 8)),
	2719 => std_logic_vector(to_unsigned(42, 8)),
	2720 => std_logic_vector(to_unsigned(42, 8)),
	2721 => std_logic_vector(to_unsigned(41, 8)),
	2722 => std_logic_vector(to_unsigned(41, 8)),
	2723 => std_logic_vector(to_unsigned(42, 8)),
	2724 => std_logic_vector(to_unsigned(42, 8)),
	2725 => std_logic_vector(to_unsigned(42, 8)),
	2726 => std_logic_vector(to_unsigned(42, 8)),
	2727 => std_logic_vector(to_unsigned(41, 8)),
	2728 => std_logic_vector(to_unsigned(41, 8)),
	2729 => std_logic_vector(to_unsigned(42, 8)),
	2730 => std_logic_vector(to_unsigned(42, 8)),
	2731 => std_logic_vector(to_unsigned(42, 8)),
	2732 => std_logic_vector(to_unsigned(41, 8)),
	2733 => std_logic_vector(to_unsigned(42, 8)),
	2734 => std_logic_vector(to_unsigned(42, 8)),
	2735 => std_logic_vector(to_unsigned(41, 8)),
	2736 => std_logic_vector(to_unsigned(42, 8)),
	2737 => std_logic_vector(to_unsigned(42, 8)),
	2738 => std_logic_vector(to_unsigned(42, 8)),
	2739 => std_logic_vector(to_unsigned(42, 8)),
	2740 => std_logic_vector(to_unsigned(42, 8)),
	2741 => std_logic_vector(to_unsigned(41, 8)),
	2742 => std_logic_vector(to_unsigned(42, 8)),
	2743 => std_logic_vector(to_unsigned(42, 8)),
	2744 => std_logic_vector(to_unsigned(41, 8)),
	2745 => std_logic_vector(to_unsigned(41, 8)),
	2746 => std_logic_vector(to_unsigned(42, 8)),
	2747 => std_logic_vector(to_unsigned(41, 8)),
	2748 => std_logic_vector(to_unsigned(41, 8)),
	2749 => std_logic_vector(to_unsigned(41, 8)),
	2750 => std_logic_vector(to_unsigned(42, 8)),
	2751 => std_logic_vector(to_unsigned(41, 8)),
	2752 => std_logic_vector(to_unsigned(41, 8)),
	2753 => std_logic_vector(to_unsigned(41, 8)),
	2754 => std_logic_vector(to_unsigned(42, 8)),
	2755 => std_logic_vector(to_unsigned(42, 8)),
	2756 => std_logic_vector(to_unsigned(42, 8)),
	2757 => std_logic_vector(to_unsigned(42, 8)),
	2758 => std_logic_vector(to_unsigned(42, 8)),
	2759 => std_logic_vector(to_unsigned(42, 8)),
	2760 => std_logic_vector(to_unsigned(42, 8)),
	2761 => std_logic_vector(to_unsigned(41, 8)),
	2762 => std_logic_vector(to_unsigned(42, 8)),
	2763 => std_logic_vector(to_unsigned(41, 8)),
	2764 => std_logic_vector(to_unsigned(42, 8)),
	2765 => std_logic_vector(to_unsigned(41, 8)),
	2766 => std_logic_vector(to_unsigned(41, 8)),
	2767 => std_logic_vector(to_unsigned(41, 8)),
	2768 => std_logic_vector(to_unsigned(42, 8)),
	2769 => std_logic_vector(to_unsigned(41, 8)),
	2770 => std_logic_vector(to_unsigned(41, 8)),
	2771 => std_logic_vector(to_unsigned(41, 8)),
	2772 => std_logic_vector(to_unsigned(42, 8)),
	2773 => std_logic_vector(to_unsigned(41, 8)),
	2774 => std_logic_vector(to_unsigned(42, 8)),
	2775 => std_logic_vector(to_unsigned(41, 8)),
	2776 => std_logic_vector(to_unsigned(42, 8)),
	2777 => std_logic_vector(to_unsigned(42, 8)),
	2778 => std_logic_vector(to_unsigned(42, 8)),
	2779 => std_logic_vector(to_unsigned(41, 8)),
	2780 => std_logic_vector(to_unsigned(41, 8)),
	2781 => std_logic_vector(to_unsigned(42, 8)),
	2782 => std_logic_vector(to_unsigned(41, 8)),
	2783 => std_logic_vector(to_unsigned(41, 8)),
	2784 => std_logic_vector(to_unsigned(41, 8)),
	2785 => std_logic_vector(to_unsigned(41, 8)),
	2786 => std_logic_vector(to_unsigned(41, 8)),
	2787 => std_logic_vector(to_unsigned(42, 8)),
	2788 => std_logic_vector(to_unsigned(41, 8)),
	2789 => std_logic_vector(to_unsigned(41, 8)),
	2790 => std_logic_vector(to_unsigned(41, 8)),
	2791 => std_logic_vector(to_unsigned(41, 8)),
	2792 => std_logic_vector(to_unsigned(42, 8)),
	2793 => std_logic_vector(to_unsigned(41, 8)),
	2794 => std_logic_vector(to_unsigned(42, 8)),
	2795 => std_logic_vector(to_unsigned(41, 8)),
	2796 => std_logic_vector(to_unsigned(42, 8)),
	2797 => std_logic_vector(to_unsigned(41, 8)),
	2798 => std_logic_vector(to_unsigned(41, 8)),
	2799 => std_logic_vector(to_unsigned(41, 8)),
	2800 => std_logic_vector(to_unsigned(41, 8)),
	2801 => std_logic_vector(to_unsigned(42, 8)),
	2802 => std_logic_vector(to_unsigned(41, 8)),
	2803 => std_logic_vector(to_unsigned(42, 8)),
	2804 => std_logic_vector(to_unsigned(42, 8)),
	2805 => std_logic_vector(to_unsigned(41, 8)),
	2806 => std_logic_vector(to_unsigned(41, 8)),
	2807 => std_logic_vector(to_unsigned(41, 8)),
	2808 => std_logic_vector(to_unsigned(42, 8)),
	2809 => std_logic_vector(to_unsigned(41, 8)),
	2810 => std_logic_vector(to_unsigned(41, 8)),
	2811 => std_logic_vector(to_unsigned(42, 8)),
	2812 => std_logic_vector(to_unsigned(42, 8)),
	2813 => std_logic_vector(to_unsigned(42, 8)),
	2814 => std_logic_vector(to_unsigned(42, 8)),
	2815 => std_logic_vector(to_unsigned(42, 8)),
	2816 => std_logic_vector(to_unsigned(42, 8)),
	2817 => std_logic_vector(to_unsigned(41, 8)),
	2818 => std_logic_vector(to_unsigned(42, 8)),
	2819 => std_logic_vector(to_unsigned(41, 8)),
	2820 => std_logic_vector(to_unsigned(41, 8)),
	2821 => std_logic_vector(to_unsigned(42, 8)),
	2822 => std_logic_vector(to_unsigned(42, 8)),
	2823 => std_logic_vector(to_unsigned(41, 8)),
	2824 => std_logic_vector(to_unsigned(42, 8)),
	2825 => std_logic_vector(to_unsigned(42, 8)),
	2826 => std_logic_vector(to_unsigned(41, 8)),
	2827 => std_logic_vector(to_unsigned(41, 8)),
	2828 => std_logic_vector(to_unsigned(42, 8)),
	2829 => std_logic_vector(to_unsigned(41, 8)),
	2830 => std_logic_vector(to_unsigned(41, 8)),
	2831 => std_logic_vector(to_unsigned(42, 8)),
	2832 => std_logic_vector(to_unsigned(42, 8)),
	2833 => std_logic_vector(to_unsigned(41, 8)),
	2834 => std_logic_vector(to_unsigned(41, 8)),
	2835 => std_logic_vector(to_unsigned(42, 8)),
	2836 => std_logic_vector(to_unsigned(41, 8)),
	2837 => std_logic_vector(to_unsigned(41, 8)),
	2838 => std_logic_vector(to_unsigned(41, 8)),
	2839 => std_logic_vector(to_unsigned(41, 8)),
	2840 => std_logic_vector(to_unsigned(41, 8)),
	2841 => std_logic_vector(to_unsigned(41, 8)),
	2842 => std_logic_vector(to_unsigned(41, 8)),
	2843 => std_logic_vector(to_unsigned(42, 8)),
	2844 => std_logic_vector(to_unsigned(41, 8)),
	2845 => std_logic_vector(to_unsigned(42, 8)),
	2846 => std_logic_vector(to_unsigned(42, 8)),
	2847 => std_logic_vector(to_unsigned(41, 8)),
	2848 => std_logic_vector(to_unsigned(41, 8)),
	2849 => std_logic_vector(to_unsigned(42, 8)),
	2850 => std_logic_vector(to_unsigned(42, 8)),
	2851 => std_logic_vector(to_unsigned(42, 8)),
	2852 => std_logic_vector(to_unsigned(42, 8)),
	2853 => std_logic_vector(to_unsigned(41, 8)),
	2854 => std_logic_vector(to_unsigned(41, 8)),
	2855 => std_logic_vector(to_unsigned(42, 8)),
	2856 => std_logic_vector(to_unsigned(42, 8)),
	2857 => std_logic_vector(to_unsigned(42, 8)),
	2858 => std_logic_vector(to_unsigned(42, 8)),
	2859 => std_logic_vector(to_unsigned(41, 8)),
	2860 => std_logic_vector(to_unsigned(41, 8)),
	2861 => std_logic_vector(to_unsigned(42, 8)),
	2862 => std_logic_vector(to_unsigned(42, 8)),
	2863 => std_logic_vector(to_unsigned(42, 8)),
	2864 => std_logic_vector(to_unsigned(41, 8)),
	2865 => std_logic_vector(to_unsigned(42, 8)),
	2866 => std_logic_vector(to_unsigned(41, 8)),
	2867 => std_logic_vector(to_unsigned(41, 8)),
	2868 => std_logic_vector(to_unsigned(42, 8)),
	2869 => std_logic_vector(to_unsigned(41, 8)),
	2870 => std_logic_vector(to_unsigned(42, 8)),
	2871 => std_logic_vector(to_unsigned(41, 8)),
	2872 => std_logic_vector(to_unsigned(41, 8)),
	2873 => std_logic_vector(to_unsigned(42, 8)),
	2874 => std_logic_vector(to_unsigned(41, 8)),
	2875 => std_logic_vector(to_unsigned(42, 8)),
	2876 => std_logic_vector(to_unsigned(42, 8)),
	2877 => std_logic_vector(to_unsigned(41, 8)),
	2878 => std_logic_vector(to_unsigned(41, 8)),
	2879 => std_logic_vector(to_unsigned(41, 8)),
	2880 => std_logic_vector(to_unsigned(41, 8)),
	2881 => std_logic_vector(to_unsigned(41, 8)),
	2882 => std_logic_vector(to_unsigned(42, 8)),
	2883 => std_logic_vector(to_unsigned(41, 8)),
	2884 => std_logic_vector(to_unsigned(41, 8)),
	2885 => std_logic_vector(to_unsigned(42, 8)),
	2886 => std_logic_vector(to_unsigned(41, 8)),
	2887 => std_logic_vector(to_unsigned(42, 8)),
	2888 => std_logic_vector(to_unsigned(41, 8)),
	2889 => std_logic_vector(to_unsigned(42, 8)),
	2890 => std_logic_vector(to_unsigned(41, 8)),
	2891 => std_logic_vector(to_unsigned(42, 8)),
	2892 => std_logic_vector(to_unsigned(42, 8)),
	2893 => std_logic_vector(to_unsigned(42, 8)),
	2894 => std_logic_vector(to_unsigned(42, 8)),
	2895 => std_logic_vector(to_unsigned(42, 8)),
	2896 => std_logic_vector(to_unsigned(42, 8)),
	2897 => std_logic_vector(to_unsigned(42, 8)),
	2898 => std_logic_vector(to_unsigned(42, 8)),
	2899 => std_logic_vector(to_unsigned(41, 8)),
	2900 => std_logic_vector(to_unsigned(41, 8)),
	2901 => std_logic_vector(to_unsigned(42, 8)),
	2902 => std_logic_vector(to_unsigned(42, 8)),
	2903 => std_logic_vector(to_unsigned(42, 8)),
	2904 => std_logic_vector(to_unsigned(41, 8)),
	2905 => std_logic_vector(to_unsigned(42, 8)),
	2906 => std_logic_vector(to_unsigned(42, 8)),
	2907 => std_logic_vector(to_unsigned(42, 8)),
	2908 => std_logic_vector(to_unsigned(42, 8)),
	2909 => std_logic_vector(to_unsigned(42, 8)),
	2910 => std_logic_vector(to_unsigned(41, 8)),
	2911 => std_logic_vector(to_unsigned(42, 8)),
	2912 => std_logic_vector(to_unsigned(42, 8)),
	2913 => std_logic_vector(to_unsigned(41, 8)),
	2914 => std_logic_vector(to_unsigned(42, 8)),
	2915 => std_logic_vector(to_unsigned(41, 8)),
	2916 => std_logic_vector(to_unsigned(42, 8)),
	2917 => std_logic_vector(to_unsigned(41, 8)),
	2918 => std_logic_vector(to_unsigned(41, 8)),
	2919 => std_logic_vector(to_unsigned(42, 8)),
	2920 => std_logic_vector(to_unsigned(41, 8)),
	2921 => std_logic_vector(to_unsigned(41, 8)),
	2922 => std_logic_vector(to_unsigned(41, 8)),
	2923 => std_logic_vector(to_unsigned(41, 8)),
	2924 => std_logic_vector(to_unsigned(42, 8)),
	2925 => std_logic_vector(to_unsigned(42, 8)),
	2926 => std_logic_vector(to_unsigned(42, 8)),
	2927 => std_logic_vector(to_unsigned(41, 8)),
	2928 => std_logic_vector(to_unsigned(42, 8)),
	2929 => std_logic_vector(to_unsigned(42, 8)),
	2930 => std_logic_vector(to_unsigned(42, 8)),
	2931 => std_logic_vector(to_unsigned(42, 8)),
	2932 => std_logic_vector(to_unsigned(42, 8)),
	2933 => std_logic_vector(to_unsigned(41, 8)),
	2934 => std_logic_vector(to_unsigned(42, 8)),
	2935 => std_logic_vector(to_unsigned(41, 8)),
	2936 => std_logic_vector(to_unsigned(41, 8)),
	2937 => std_logic_vector(to_unsigned(42, 8)),
	2938 => std_logic_vector(to_unsigned(42, 8)),
	2939 => std_logic_vector(to_unsigned(42, 8)),
	2940 => std_logic_vector(to_unsigned(41, 8)),
	2941 => std_logic_vector(to_unsigned(41, 8)),
	2942 => std_logic_vector(to_unsigned(42, 8)),
	2943 => std_logic_vector(to_unsigned(42, 8)),
	2944 => std_logic_vector(to_unsigned(41, 8)),
	2945 => std_logic_vector(to_unsigned(42, 8)),
	2946 => std_logic_vector(to_unsigned(41, 8)),
	2947 => std_logic_vector(to_unsigned(41, 8)),
	2948 => std_logic_vector(to_unsigned(41, 8)),
	2949 => std_logic_vector(to_unsigned(42, 8)),
	2950 => std_logic_vector(to_unsigned(42, 8)),
	2951 => std_logic_vector(to_unsigned(41, 8)),
	2952 => std_logic_vector(to_unsigned(41, 8)),
	2953 => std_logic_vector(to_unsigned(42, 8)),
	2954 => std_logic_vector(to_unsigned(42, 8)),
	2955 => std_logic_vector(to_unsigned(42, 8)),
	2956 => std_logic_vector(to_unsigned(42, 8)),
	2957 => std_logic_vector(to_unsigned(42, 8)),
	2958 => std_logic_vector(to_unsigned(42, 8)),
	2959 => std_logic_vector(to_unsigned(41, 8)),
	2960 => std_logic_vector(to_unsigned(42, 8)),
	2961 => std_logic_vector(to_unsigned(41, 8)),
	2962 => std_logic_vector(to_unsigned(42, 8)),
	2963 => std_logic_vector(to_unsigned(42, 8)),
	2964 => std_logic_vector(to_unsigned(42, 8)),
	2965 => std_logic_vector(to_unsigned(42, 8)),
	2966 => std_logic_vector(to_unsigned(42, 8)),
	2967 => std_logic_vector(to_unsigned(41, 8)),
	2968 => std_logic_vector(to_unsigned(42, 8)),
	2969 => std_logic_vector(to_unsigned(42, 8)),
	2970 => std_logic_vector(to_unsigned(41, 8)),
	2971 => std_logic_vector(to_unsigned(41, 8)),
	2972 => std_logic_vector(to_unsigned(42, 8)),
	2973 => std_logic_vector(to_unsigned(41, 8)),
	2974 => std_logic_vector(to_unsigned(41, 8)),
	2975 => std_logic_vector(to_unsigned(42, 8)),
	2976 => std_logic_vector(to_unsigned(41, 8)),
	2977 => std_logic_vector(to_unsigned(42, 8)),
	2978 => std_logic_vector(to_unsigned(42, 8)),
	2979 => std_logic_vector(to_unsigned(42, 8)),
	2980 => std_logic_vector(to_unsigned(42, 8)),
	2981 => std_logic_vector(to_unsigned(42, 8)),
	2982 => std_logic_vector(to_unsigned(42, 8)),
	2983 => std_logic_vector(to_unsigned(42, 8)),
	2984 => std_logic_vector(to_unsigned(42, 8)),
	2985 => std_logic_vector(to_unsigned(42, 8)),
	2986 => std_logic_vector(to_unsigned(41, 8)),
	2987 => std_logic_vector(to_unsigned(41, 8)),
	2988 => std_logic_vector(to_unsigned(42, 8)),
	2989 => std_logic_vector(to_unsigned(41, 8)),
	2990 => std_logic_vector(to_unsigned(41, 8)),
	2991 => std_logic_vector(to_unsigned(41, 8)),
	2992 => std_logic_vector(to_unsigned(41, 8)),
	2993 => std_logic_vector(to_unsigned(42, 8)),
	2994 => std_logic_vector(to_unsigned(42, 8)),
	2995 => std_logic_vector(to_unsigned(41, 8)),
	2996 => std_logic_vector(to_unsigned(42, 8)),
	2997 => std_logic_vector(to_unsigned(41, 8)),
	2998 => std_logic_vector(to_unsigned(42, 8)),
	2999 => std_logic_vector(to_unsigned(42, 8)),
	3000 => std_logic_vector(to_unsigned(42, 8)),
	3001 => std_logic_vector(to_unsigned(42, 8)),
	3002 => std_logic_vector(to_unsigned(42, 8)),
	3003 => std_logic_vector(to_unsigned(41, 8)),
	3004 => std_logic_vector(to_unsigned(41, 8)),
	3005 => std_logic_vector(to_unsigned(41, 8)),
	3006 => std_logic_vector(to_unsigned(41, 8)),
	3007 => std_logic_vector(to_unsigned(42, 8)),
	3008 => std_logic_vector(to_unsigned(41, 8)),
	3009 => std_logic_vector(to_unsigned(41, 8)),
	3010 => std_logic_vector(to_unsigned(41, 8)),
	3011 => std_logic_vector(to_unsigned(42, 8)),
	3012 => std_logic_vector(to_unsigned(42, 8)),
	3013 => std_logic_vector(to_unsigned(42, 8)),
	3014 => std_logic_vector(to_unsigned(42, 8)),
	3015 => std_logic_vector(to_unsigned(42, 8)),
	3016 => std_logic_vector(to_unsigned(42, 8)),
	3017 => std_logic_vector(to_unsigned(42, 8)),
	3018 => std_logic_vector(to_unsigned(42, 8)),
	3019 => std_logic_vector(to_unsigned(42, 8)),
	3020 => std_logic_vector(to_unsigned(42, 8)),
	3021 => std_logic_vector(to_unsigned(41, 8)),
	3022 => std_logic_vector(to_unsigned(41, 8)),
	3023 => std_logic_vector(to_unsigned(41, 8)),
	3024 => std_logic_vector(to_unsigned(42, 8)),
	3025 => std_logic_vector(to_unsigned(41, 8)),
	3026 => std_logic_vector(to_unsigned(42, 8)),
	3027 => std_logic_vector(to_unsigned(41, 8)),
	3028 => std_logic_vector(to_unsigned(41, 8)),
	3029 => std_logic_vector(to_unsigned(41, 8)),
	3030 => std_logic_vector(to_unsigned(41, 8)),
	3031 => std_logic_vector(to_unsigned(41, 8)),
	3032 => std_logic_vector(to_unsigned(41, 8)),
	3033 => std_logic_vector(to_unsigned(42, 8)),
	3034 => std_logic_vector(to_unsigned(42, 8)),
	3035 => std_logic_vector(to_unsigned(41, 8)),
	3036 => std_logic_vector(to_unsigned(41, 8)),
	3037 => std_logic_vector(to_unsigned(42, 8)),
	3038 => std_logic_vector(to_unsigned(42, 8)),
	3039 => std_logic_vector(to_unsigned(41, 8)),
	3040 => std_logic_vector(to_unsigned(41, 8)),
	3041 => std_logic_vector(to_unsigned(41, 8)),
	3042 => std_logic_vector(to_unsigned(42, 8)),
	3043 => std_logic_vector(to_unsigned(42, 8)),
	3044 => std_logic_vector(to_unsigned(41, 8)),
	3045 => std_logic_vector(to_unsigned(41, 8)),
	3046 => std_logic_vector(to_unsigned(42, 8)),
	3047 => std_logic_vector(to_unsigned(42, 8)),
	3048 => std_logic_vector(to_unsigned(41, 8)),
	3049 => std_logic_vector(to_unsigned(42, 8)),
	3050 => std_logic_vector(to_unsigned(42, 8)),
	3051 => std_logic_vector(to_unsigned(41, 8)),
	3052 => std_logic_vector(to_unsigned(41, 8)),
	3053 => std_logic_vector(to_unsigned(42, 8)),
	3054 => std_logic_vector(to_unsigned(42, 8)),
	3055 => std_logic_vector(to_unsigned(41, 8)),
	3056 => std_logic_vector(to_unsigned(42, 8)),
	3057 => std_logic_vector(to_unsigned(41, 8)),
	3058 => std_logic_vector(to_unsigned(42, 8)),
	3059 => std_logic_vector(to_unsigned(42, 8)),
	3060 => std_logic_vector(to_unsigned(42, 8)),
	3061 => std_logic_vector(to_unsigned(41, 8)),
	3062 => std_logic_vector(to_unsigned(41, 8)),
	3063 => std_logic_vector(to_unsigned(42, 8)),
	3064 => std_logic_vector(to_unsigned(42, 8)),
	3065 => std_logic_vector(to_unsigned(41, 8)),
	3066 => std_logic_vector(to_unsigned(41, 8)),
	3067 => std_logic_vector(to_unsigned(41, 8)),
	3068 => std_logic_vector(to_unsigned(41, 8)),
	3069 => std_logic_vector(to_unsigned(41, 8)),
	3070 => std_logic_vector(to_unsigned(42, 8)),
	3071 => std_logic_vector(to_unsigned(42, 8)),
	3072 => std_logic_vector(to_unsigned(42, 8)),
	3073 => std_logic_vector(to_unsigned(41, 8)),
	3074 => std_logic_vector(to_unsigned(41, 8)),
	3075 => std_logic_vector(to_unsigned(41, 8)),
	3076 => std_logic_vector(to_unsigned(42, 8)),
	3077 => std_logic_vector(to_unsigned(42, 8)),
	3078 => std_logic_vector(to_unsigned(41, 8)),
	3079 => std_logic_vector(to_unsigned(41, 8)),
	3080 => std_logic_vector(to_unsigned(42, 8)),
	3081 => std_logic_vector(to_unsigned(41, 8)),
	3082 => std_logic_vector(to_unsigned(41, 8)),
	3083 => std_logic_vector(to_unsigned(41, 8)),
	3084 => std_logic_vector(to_unsigned(42, 8)),
	3085 => std_logic_vector(to_unsigned(41, 8)),
	3086 => std_logic_vector(to_unsigned(41, 8)),
	3087 => std_logic_vector(to_unsigned(42, 8)),
	3088 => std_logic_vector(to_unsigned(42, 8)),
	3089 => std_logic_vector(to_unsigned(42, 8)),
	3090 => std_logic_vector(to_unsigned(41, 8)),
	3091 => std_logic_vector(to_unsigned(42, 8)),
	3092 => std_logic_vector(to_unsigned(41, 8)),
	3093 => std_logic_vector(to_unsigned(41, 8)),
	3094 => std_logic_vector(to_unsigned(42, 8)),
	3095 => std_logic_vector(to_unsigned(41, 8)),
	3096 => std_logic_vector(to_unsigned(41, 8)),
	3097 => std_logic_vector(to_unsigned(42, 8)),
	3098 => std_logic_vector(to_unsigned(41, 8)),
	3099 => std_logic_vector(to_unsigned(42, 8)),
	3100 => std_logic_vector(to_unsigned(42, 8)),
	3101 => std_logic_vector(to_unsigned(42, 8)),
	3102 => std_logic_vector(to_unsigned(42, 8)),
	3103 => std_logic_vector(to_unsigned(41, 8)),
	3104 => std_logic_vector(to_unsigned(42, 8)),
	3105 => std_logic_vector(to_unsigned(42, 8)),
	3106 => std_logic_vector(to_unsigned(41, 8)),
	3107 => std_logic_vector(to_unsigned(42, 8)),
	3108 => std_logic_vector(to_unsigned(41, 8)),
	3109 => std_logic_vector(to_unsigned(42, 8)),
	3110 => std_logic_vector(to_unsigned(42, 8)),
	3111 => std_logic_vector(to_unsigned(41, 8)),
	3112 => std_logic_vector(to_unsigned(41, 8)),
	3113 => std_logic_vector(to_unsigned(41, 8)),
	3114 => std_logic_vector(to_unsigned(42, 8)),
	3115 => std_logic_vector(to_unsigned(42, 8)),
	3116 => std_logic_vector(to_unsigned(41, 8)),
	3117 => std_logic_vector(to_unsigned(41, 8)),
	3118 => std_logic_vector(to_unsigned(41, 8)),
	3119 => std_logic_vector(to_unsigned(42, 8)),
	3120 => std_logic_vector(to_unsigned(42, 8)),
	3121 => std_logic_vector(to_unsigned(42, 8)),
	3122 => std_logic_vector(to_unsigned(42, 8)),
	3123 => std_logic_vector(to_unsigned(41, 8)),
	3124 => std_logic_vector(to_unsigned(42, 8)),
	3125 => std_logic_vector(to_unsigned(41, 8)),
	3126 => std_logic_vector(to_unsigned(41, 8)),
	3127 => std_logic_vector(to_unsigned(42, 8)),
	3128 => std_logic_vector(to_unsigned(41, 8)),
	3129 => std_logic_vector(to_unsigned(41, 8)),
	3130 => std_logic_vector(to_unsigned(41, 8)),
	3131 => std_logic_vector(to_unsigned(42, 8)),
	3132 => std_logic_vector(to_unsigned(42, 8)),
	3133 => std_logic_vector(to_unsigned(41, 8)),
	3134 => std_logic_vector(to_unsigned(41, 8)),
	3135 => std_logic_vector(to_unsigned(42, 8)),
	3136 => std_logic_vector(to_unsigned(41, 8)),
	3137 => std_logic_vector(to_unsigned(42, 8)),
	3138 => std_logic_vector(to_unsigned(42, 8)),
	3139 => std_logic_vector(to_unsigned(41, 8)),
	3140 => std_logic_vector(to_unsigned(42, 8)),
	3141 => std_logic_vector(to_unsigned(42, 8)),
	3142 => std_logic_vector(to_unsigned(42, 8)),
	3143 => std_logic_vector(to_unsigned(42, 8)),
	3144 => std_logic_vector(to_unsigned(41, 8)),
	3145 => std_logic_vector(to_unsigned(42, 8)),
	3146 => std_logic_vector(to_unsigned(42, 8)),
	3147 => std_logic_vector(to_unsigned(42, 8)),
	3148 => std_logic_vector(to_unsigned(41, 8)),
	3149 => std_logic_vector(to_unsigned(42, 8)),
	3150 => std_logic_vector(to_unsigned(41, 8)),
	3151 => std_logic_vector(to_unsigned(41, 8)),
	3152 => std_logic_vector(to_unsigned(41, 8)),
	3153 => std_logic_vector(to_unsigned(41, 8)),
	3154 => std_logic_vector(to_unsigned(41, 8)),
	3155 => std_logic_vector(to_unsigned(41, 8)),
	3156 => std_logic_vector(to_unsigned(41, 8)),
	3157 => std_logic_vector(to_unsigned(42, 8)),
	3158 => std_logic_vector(to_unsigned(42, 8)),
	3159 => std_logic_vector(to_unsigned(42, 8)),
	3160 => std_logic_vector(to_unsigned(42, 8)),
	3161 => std_logic_vector(to_unsigned(42, 8)),
	3162 => std_logic_vector(to_unsigned(42, 8)),
	3163 => std_logic_vector(to_unsigned(42, 8)),
	3164 => std_logic_vector(to_unsigned(41, 8)),
	3165 => std_logic_vector(to_unsigned(41, 8)),
	3166 => std_logic_vector(to_unsigned(41, 8)),
	3167 => std_logic_vector(to_unsigned(41, 8)),
	3168 => std_logic_vector(to_unsigned(41, 8)),
	3169 => std_logic_vector(to_unsigned(42, 8)),
	3170 => std_logic_vector(to_unsigned(41, 8)),
	3171 => std_logic_vector(to_unsigned(42, 8)),
	3172 => std_logic_vector(to_unsigned(41, 8)),
	3173 => std_logic_vector(to_unsigned(42, 8)),
	3174 => std_logic_vector(to_unsigned(41, 8)),
	3175 => std_logic_vector(to_unsigned(42, 8)),
	3176 => std_logic_vector(to_unsigned(42, 8)),
	3177 => std_logic_vector(to_unsigned(41, 8)),
	3178 => std_logic_vector(to_unsigned(41, 8)),
	3179 => std_logic_vector(to_unsigned(42, 8)),
	3180 => std_logic_vector(to_unsigned(41, 8)),
	3181 => std_logic_vector(to_unsigned(41, 8)),
	3182 => std_logic_vector(to_unsigned(42, 8)),
	3183 => std_logic_vector(to_unsigned(42, 8)),
	3184 => std_logic_vector(to_unsigned(42, 8)),
	3185 => std_logic_vector(to_unsigned(42, 8)),
	3186 => std_logic_vector(to_unsigned(42, 8)),
	3187 => std_logic_vector(to_unsigned(42, 8)),
	3188 => std_logic_vector(to_unsigned(42, 8)),
	3189 => std_logic_vector(to_unsigned(42, 8)),
	3190 => std_logic_vector(to_unsigned(42, 8)),
	3191 => std_logic_vector(to_unsigned(41, 8)),
	3192 => std_logic_vector(to_unsigned(41, 8)),
	3193 => std_logic_vector(to_unsigned(42, 8)),
	3194 => std_logic_vector(to_unsigned(41, 8)),
	3195 => std_logic_vector(to_unsigned(42, 8)),
	3196 => std_logic_vector(to_unsigned(42, 8)),
	3197 => std_logic_vector(to_unsigned(41, 8)),
	3198 => std_logic_vector(to_unsigned(42, 8)),
	3199 => std_logic_vector(to_unsigned(41, 8)),
	3200 => std_logic_vector(to_unsigned(41, 8)),
	3201 => std_logic_vector(to_unsigned(41, 8)),
	3202 => std_logic_vector(to_unsigned(42, 8)),
	3203 => std_logic_vector(to_unsigned(42, 8)),
	3204 => std_logic_vector(to_unsigned(42, 8)),
	3205 => std_logic_vector(to_unsigned(41, 8)),
	3206 => std_logic_vector(to_unsigned(41, 8)),
	3207 => std_logic_vector(to_unsigned(41, 8)),
	3208 => std_logic_vector(to_unsigned(41, 8)),
	3209 => std_logic_vector(to_unsigned(41, 8)),
	3210 => std_logic_vector(to_unsigned(42, 8)),
	3211 => std_logic_vector(to_unsigned(42, 8)),
	3212 => std_logic_vector(to_unsigned(41, 8)),
	3213 => std_logic_vector(to_unsigned(41, 8)),
	3214 => std_logic_vector(to_unsigned(41, 8)),
	3215 => std_logic_vector(to_unsigned(42, 8)),
	3216 => std_logic_vector(to_unsigned(41, 8)),
	3217 => std_logic_vector(to_unsigned(42, 8)),
	3218 => std_logic_vector(to_unsigned(41, 8)),
	3219 => std_logic_vector(to_unsigned(42, 8)),
	3220 => std_logic_vector(to_unsigned(41, 8)),
	3221 => std_logic_vector(to_unsigned(41, 8)),
	3222 => std_logic_vector(to_unsigned(42, 8)),
	3223 => std_logic_vector(to_unsigned(42, 8)),
	3224 => std_logic_vector(to_unsigned(41, 8)),
	3225 => std_logic_vector(to_unsigned(41, 8)),
	3226 => std_logic_vector(to_unsigned(42, 8)),
	3227 => std_logic_vector(to_unsigned(42, 8)),
	3228 => std_logic_vector(to_unsigned(42, 8)),
	3229 => std_logic_vector(to_unsigned(41, 8)),
	3230 => std_logic_vector(to_unsigned(41, 8)),
	3231 => std_logic_vector(to_unsigned(41, 8)),
	3232 => std_logic_vector(to_unsigned(42, 8)),
	3233 => std_logic_vector(to_unsigned(42, 8)),
	3234 => std_logic_vector(to_unsigned(41, 8)),
	3235 => std_logic_vector(to_unsigned(42, 8)),
	3236 => std_logic_vector(to_unsigned(41, 8)),
	3237 => std_logic_vector(to_unsigned(42, 8)),
	3238 => std_logic_vector(to_unsigned(42, 8)),
	3239 => std_logic_vector(to_unsigned(42, 8)),
	3240 => std_logic_vector(to_unsigned(41, 8)),
	3241 => std_logic_vector(to_unsigned(41, 8)),
	3242 => std_logic_vector(to_unsigned(41, 8)),
	3243 => std_logic_vector(to_unsigned(41, 8)),
	3244 => std_logic_vector(to_unsigned(41, 8)),
	3245 => std_logic_vector(to_unsigned(41, 8)),
	3246 => std_logic_vector(to_unsigned(41, 8)),
	3247 => std_logic_vector(to_unsigned(42, 8)),
	3248 => std_logic_vector(to_unsigned(41, 8)),
	3249 => std_logic_vector(to_unsigned(42, 8)),
	3250 => std_logic_vector(to_unsigned(42, 8)),
	3251 => std_logic_vector(to_unsigned(42, 8)),
	3252 => std_logic_vector(to_unsigned(42, 8)),
	3253 => std_logic_vector(to_unsigned(42, 8)),
	3254 => std_logic_vector(to_unsigned(42, 8)),
	3255 => std_logic_vector(to_unsigned(41, 8)),
	3256 => std_logic_vector(to_unsigned(41, 8)),
	3257 => std_logic_vector(to_unsigned(42, 8)),
	3258 => std_logic_vector(to_unsigned(41, 8)),
	3259 => std_logic_vector(to_unsigned(41, 8)),
	3260 => std_logic_vector(to_unsigned(42, 8)),
	3261 => std_logic_vector(to_unsigned(41, 8)),
	3262 => std_logic_vector(to_unsigned(41, 8)),
	3263 => std_logic_vector(to_unsigned(41, 8)),
	3264 => std_logic_vector(to_unsigned(41, 8)),
	3265 => std_logic_vector(to_unsigned(41, 8)),
	3266 => std_logic_vector(to_unsigned(41, 8)),
	3267 => std_logic_vector(to_unsigned(41, 8)),
	3268 => std_logic_vector(to_unsigned(41, 8)),
	3269 => std_logic_vector(to_unsigned(42, 8)),
	3270 => std_logic_vector(to_unsigned(41, 8)),
	3271 => std_logic_vector(to_unsigned(41, 8)),
	3272 => std_logic_vector(to_unsigned(42, 8)),
	3273 => std_logic_vector(to_unsigned(41, 8)),
	3274 => std_logic_vector(to_unsigned(41, 8)),
	3275 => std_logic_vector(to_unsigned(42, 8)),
	3276 => std_logic_vector(to_unsigned(41, 8)),
	3277 => std_logic_vector(to_unsigned(41, 8)),
	3278 => std_logic_vector(to_unsigned(41, 8)),
	3279 => std_logic_vector(to_unsigned(41, 8)),
	3280 => std_logic_vector(to_unsigned(42, 8)),
	3281 => std_logic_vector(to_unsigned(41, 8)),
	3282 => std_logic_vector(to_unsigned(42, 8)),
	3283 => std_logic_vector(to_unsigned(41, 8)),
	3284 => std_logic_vector(to_unsigned(42, 8)),
	3285 => std_logic_vector(to_unsigned(41, 8)),
	3286 => std_logic_vector(to_unsigned(41, 8)),
	3287 => std_logic_vector(to_unsigned(41, 8)),
	3288 => std_logic_vector(to_unsigned(42, 8)),
	3289 => std_logic_vector(to_unsigned(42, 8)),
	3290 => std_logic_vector(to_unsigned(41, 8)),
	3291 => std_logic_vector(to_unsigned(42, 8)),
	3292 => std_logic_vector(to_unsigned(41, 8)),
	3293 => std_logic_vector(to_unsigned(41, 8)),
	3294 => std_logic_vector(to_unsigned(42, 8)),
	3295 => std_logic_vector(to_unsigned(41, 8)),
	3296 => std_logic_vector(to_unsigned(41, 8)),
	3297 => std_logic_vector(to_unsigned(42, 8)),
	3298 => std_logic_vector(to_unsigned(41, 8)),
	3299 => std_logic_vector(to_unsigned(41, 8)),
	3300 => std_logic_vector(to_unsigned(42, 8)),
	3301 => std_logic_vector(to_unsigned(42, 8)),
	3302 => std_logic_vector(to_unsigned(42, 8)),
	3303 => std_logic_vector(to_unsigned(42, 8)),
	3304 => std_logic_vector(to_unsigned(41, 8)),
	3305 => std_logic_vector(to_unsigned(42, 8)),
	3306 => std_logic_vector(to_unsigned(41, 8)),
	3307 => std_logic_vector(to_unsigned(41, 8)),
	3308 => std_logic_vector(to_unsigned(41, 8)),
	3309 => std_logic_vector(to_unsigned(41, 8)),
	3310 => std_logic_vector(to_unsigned(41, 8)),
	3311 => std_logic_vector(to_unsigned(42, 8)),
	3312 => std_logic_vector(to_unsigned(41, 8)),
	3313 => std_logic_vector(to_unsigned(41, 8)),
	3314 => std_logic_vector(to_unsigned(42, 8)),
	3315 => std_logic_vector(to_unsigned(41, 8)),
	3316 => std_logic_vector(to_unsigned(42, 8)),
	3317 => std_logic_vector(to_unsigned(42, 8)),
	3318 => std_logic_vector(to_unsigned(42, 8)),
	3319 => std_logic_vector(to_unsigned(42, 8)),
	3320 => std_logic_vector(to_unsigned(41, 8)),
	3321 => std_logic_vector(to_unsigned(41, 8)),
	3322 => std_logic_vector(to_unsigned(42, 8)),
	3323 => std_logic_vector(to_unsigned(41, 8)),
	3324 => std_logic_vector(to_unsigned(42, 8)),
	3325 => std_logic_vector(to_unsigned(42, 8)),
	3326 => std_logic_vector(to_unsigned(42, 8)),
	3327 => std_logic_vector(to_unsigned(41, 8)),
	3328 => std_logic_vector(to_unsigned(41, 8)),
	3329 => std_logic_vector(to_unsigned(42, 8)),
	3330 => std_logic_vector(to_unsigned(42, 8)),
	3331 => std_logic_vector(to_unsigned(42, 8)),
	3332 => std_logic_vector(to_unsigned(41, 8)),
	3333 => std_logic_vector(to_unsigned(42, 8)),
	3334 => std_logic_vector(to_unsigned(42, 8)),
	3335 => std_logic_vector(to_unsigned(42, 8)),
	3336 => std_logic_vector(to_unsigned(41, 8)),
	3337 => std_logic_vector(to_unsigned(41, 8)),
	3338 => std_logic_vector(to_unsigned(42, 8)),
	3339 => std_logic_vector(to_unsigned(42, 8)),
	3340 => std_logic_vector(to_unsigned(41, 8)),
	3341 => std_logic_vector(to_unsigned(41, 8)),
	3342 => std_logic_vector(to_unsigned(42, 8)),
	3343 => std_logic_vector(to_unsigned(42, 8)),
	3344 => std_logic_vector(to_unsigned(42, 8)),
	3345 => std_logic_vector(to_unsigned(42, 8)),
	3346 => std_logic_vector(to_unsigned(41, 8)),
	3347 => std_logic_vector(to_unsigned(41, 8)),
	3348 => std_logic_vector(to_unsigned(42, 8)),
	3349 => std_logic_vector(to_unsigned(41, 8)),
	3350 => std_logic_vector(to_unsigned(42, 8)),
	3351 => std_logic_vector(to_unsigned(41, 8)),
	3352 => std_logic_vector(to_unsigned(41, 8)),
	3353 => std_logic_vector(to_unsigned(42, 8)),
	3354 => std_logic_vector(to_unsigned(41, 8)),
	3355 => std_logic_vector(to_unsigned(42, 8)),
	3356 => std_logic_vector(to_unsigned(42, 8)),
	3357 => std_logic_vector(to_unsigned(41, 8)),
	3358 => std_logic_vector(to_unsigned(41, 8)),
	3359 => std_logic_vector(to_unsigned(42, 8)),
	3360 => std_logic_vector(to_unsigned(42, 8)),
	3361 => std_logic_vector(to_unsigned(41, 8)),
	3362 => std_logic_vector(to_unsigned(42, 8)),
	3363 => std_logic_vector(to_unsigned(41, 8)),
	3364 => std_logic_vector(to_unsigned(41, 8)),
	3365 => std_logic_vector(to_unsigned(41, 8)),
	3366 => std_logic_vector(to_unsigned(41, 8)),
	3367 => std_logic_vector(to_unsigned(42, 8)),
	3368 => std_logic_vector(to_unsigned(42, 8)),
	3369 => std_logic_vector(to_unsigned(41, 8)),
	3370 => std_logic_vector(to_unsigned(41, 8)),
	3371 => std_logic_vector(to_unsigned(41, 8)),
	3372 => std_logic_vector(to_unsigned(41, 8)),
	3373 => std_logic_vector(to_unsigned(41, 8)),
	3374 => std_logic_vector(to_unsigned(42, 8)),
	3375 => std_logic_vector(to_unsigned(42, 8)),
	3376 => std_logic_vector(to_unsigned(42, 8)),
	3377 => std_logic_vector(to_unsigned(41, 8)),
	3378 => std_logic_vector(to_unsigned(41, 8)),
	3379 => std_logic_vector(to_unsigned(41, 8)),
	3380 => std_logic_vector(to_unsigned(42, 8)),
	3381 => std_logic_vector(to_unsigned(42, 8)),
	3382 => std_logic_vector(to_unsigned(42, 8)),
	3383 => std_logic_vector(to_unsigned(42, 8)),
	3384 => std_logic_vector(to_unsigned(42, 8)),
	3385 => std_logic_vector(to_unsigned(42, 8)),
	3386 => std_logic_vector(to_unsigned(42, 8)),
	3387 => std_logic_vector(to_unsigned(42, 8)),
	3388 => std_logic_vector(to_unsigned(41, 8)),
	3389 => std_logic_vector(to_unsigned(42, 8)),
	3390 => std_logic_vector(to_unsigned(41, 8)),
	3391 => std_logic_vector(to_unsigned(42, 8)),
	3392 => std_logic_vector(to_unsigned(42, 8)),
	3393 => std_logic_vector(to_unsigned(41, 8)),
	3394 => std_logic_vector(to_unsigned(41, 8)),
	3395 => std_logic_vector(to_unsigned(41, 8)),
	3396 => std_logic_vector(to_unsigned(41, 8)),
	3397 => std_logic_vector(to_unsigned(41, 8)),
	3398 => std_logic_vector(to_unsigned(42, 8)),
	3399 => std_logic_vector(to_unsigned(42, 8)),
	3400 => std_logic_vector(to_unsigned(42, 8)),
	3401 => std_logic_vector(to_unsigned(42, 8)),
	3402 => std_logic_vector(to_unsigned(41, 8)),
	3403 => std_logic_vector(to_unsigned(42, 8)),
	3404 => std_logic_vector(to_unsigned(42, 8)),
	3405 => std_logic_vector(to_unsigned(41, 8)),
	3406 => std_logic_vector(to_unsigned(41, 8)),
	3407 => std_logic_vector(to_unsigned(42, 8)),
	3408 => std_logic_vector(to_unsigned(41, 8)),
	3409 => std_logic_vector(to_unsigned(41, 8)),
	3410 => std_logic_vector(to_unsigned(41, 8)),
	3411 => std_logic_vector(to_unsigned(42, 8)),
	3412 => std_logic_vector(to_unsigned(42, 8)),
	3413 => std_logic_vector(to_unsigned(42, 8)),
	3414 => std_logic_vector(to_unsigned(42, 8)),
	3415 => std_logic_vector(to_unsigned(41, 8)),
	3416 => std_logic_vector(to_unsigned(41, 8)),
	3417 => std_logic_vector(to_unsigned(41, 8)),
	3418 => std_logic_vector(to_unsigned(42, 8)),
	3419 => std_logic_vector(to_unsigned(41, 8)),
	3420 => std_logic_vector(to_unsigned(41, 8)),
	3421 => std_logic_vector(to_unsigned(41, 8)),
	3422 => std_logic_vector(to_unsigned(41, 8)),
	3423 => std_logic_vector(to_unsigned(42, 8)),
	3424 => std_logic_vector(to_unsigned(42, 8)),
	3425 => std_logic_vector(to_unsigned(42, 8)),
	3426 => std_logic_vector(to_unsigned(42, 8)),
	3427 => std_logic_vector(to_unsigned(42, 8)),
	3428 => std_logic_vector(to_unsigned(42, 8)),
	3429 => std_logic_vector(to_unsigned(42, 8)),
	3430 => std_logic_vector(to_unsigned(41, 8)),
	3431 => std_logic_vector(to_unsigned(42, 8)),
	3432 => std_logic_vector(to_unsigned(42, 8)),
	3433 => std_logic_vector(to_unsigned(41, 8)),
	3434 => std_logic_vector(to_unsigned(42, 8)),
	3435 => std_logic_vector(to_unsigned(41, 8)),
	3436 => std_logic_vector(to_unsigned(41, 8)),
	3437 => std_logic_vector(to_unsigned(42, 8)),
	3438 => std_logic_vector(to_unsigned(41, 8)),
	3439 => std_logic_vector(to_unsigned(42, 8)),
	3440 => std_logic_vector(to_unsigned(42, 8)),
	3441 => std_logic_vector(to_unsigned(41, 8)),
	3442 => std_logic_vector(to_unsigned(41, 8)),
	3443 => std_logic_vector(to_unsigned(41, 8)),
	3444 => std_logic_vector(to_unsigned(41, 8)),
	3445 => std_logic_vector(to_unsigned(42, 8)),
	3446 => std_logic_vector(to_unsigned(42, 8)),
	3447 => std_logic_vector(to_unsigned(41, 8)),
	3448 => std_logic_vector(to_unsigned(42, 8)),
	3449 => std_logic_vector(to_unsigned(42, 8)),
	3450 => std_logic_vector(to_unsigned(41, 8)),
	3451 => std_logic_vector(to_unsigned(41, 8)),
	3452 => std_logic_vector(to_unsigned(42, 8)),
	3453 => std_logic_vector(to_unsigned(41, 8)),
	3454 => std_logic_vector(to_unsigned(42, 8)),
	3455 => std_logic_vector(to_unsigned(42, 8)),
	3456 => std_logic_vector(to_unsigned(42, 8)),
	3457 => std_logic_vector(to_unsigned(41, 8)),
	3458 => std_logic_vector(to_unsigned(42, 8)),
	3459 => std_logic_vector(to_unsigned(41, 8)),
	3460 => std_logic_vector(to_unsigned(42, 8)),
	3461 => std_logic_vector(to_unsigned(41, 8)),
	3462 => std_logic_vector(to_unsigned(41, 8)),
	3463 => std_logic_vector(to_unsigned(42, 8)),
	3464 => std_logic_vector(to_unsigned(42, 8)),
	3465 => std_logic_vector(to_unsigned(41, 8)),
	3466 => std_logic_vector(to_unsigned(42, 8)),
	3467 => std_logic_vector(to_unsigned(42, 8)),
	3468 => std_logic_vector(to_unsigned(42, 8)),
	3469 => std_logic_vector(to_unsigned(41, 8)),
	3470 => std_logic_vector(to_unsigned(41, 8)),
	3471 => std_logic_vector(to_unsigned(42, 8)),
	3472 => std_logic_vector(to_unsigned(42, 8)),
	3473 => std_logic_vector(to_unsigned(42, 8)),
	3474 => std_logic_vector(to_unsigned(42, 8)),
	3475 => std_logic_vector(to_unsigned(41, 8)),
	3476 => std_logic_vector(to_unsigned(42, 8)),
	3477 => std_logic_vector(to_unsigned(42, 8)),
	3478 => std_logic_vector(to_unsigned(41, 8)),
	3479 => std_logic_vector(to_unsigned(41, 8)),
	3480 => std_logic_vector(to_unsigned(41, 8)),
	3481 => std_logic_vector(to_unsigned(41, 8)),
	3482 => std_logic_vector(to_unsigned(42, 8)),
	3483 => std_logic_vector(to_unsigned(42, 8)),
	3484 => std_logic_vector(to_unsigned(41, 8)),
	3485 => std_logic_vector(to_unsigned(41, 8)),
	3486 => std_logic_vector(to_unsigned(42, 8)),
	3487 => std_logic_vector(to_unsigned(41, 8)),
	3488 => std_logic_vector(to_unsigned(41, 8)),
	3489 => std_logic_vector(to_unsigned(41, 8)),
	3490 => std_logic_vector(to_unsigned(41, 8)),
	3491 => std_logic_vector(to_unsigned(41, 8)),
	3492 => std_logic_vector(to_unsigned(42, 8)),
	3493 => std_logic_vector(to_unsigned(41, 8)),
	3494 => std_logic_vector(to_unsigned(41, 8)),
	3495 => std_logic_vector(to_unsigned(41, 8)),
	3496 => std_logic_vector(to_unsigned(42, 8)),
	3497 => std_logic_vector(to_unsigned(41, 8)),
	3498 => std_logic_vector(to_unsigned(41, 8)),
	3499 => std_logic_vector(to_unsigned(42, 8)),
	3500 => std_logic_vector(to_unsigned(41, 8)),
	3501 => std_logic_vector(to_unsigned(42, 8)),
	3502 => std_logic_vector(to_unsigned(41, 8)),
	3503 => std_logic_vector(to_unsigned(42, 8)),
	3504 => std_logic_vector(to_unsigned(42, 8)),
	3505 => std_logic_vector(to_unsigned(42, 8)),
	3506 => std_logic_vector(to_unsigned(41, 8)),
	3507 => std_logic_vector(to_unsigned(42, 8)),
	3508 => std_logic_vector(to_unsigned(41, 8)),
	3509 => std_logic_vector(to_unsigned(42, 8)),
	3510 => std_logic_vector(to_unsigned(41, 8)),
	3511 => std_logic_vector(to_unsigned(42, 8)),
	3512 => std_logic_vector(to_unsigned(41, 8)),
	3513 => std_logic_vector(to_unsigned(42, 8)),
	3514 => std_logic_vector(to_unsigned(42, 8)),
	3515 => std_logic_vector(to_unsigned(42, 8)),
	3516 => std_logic_vector(to_unsigned(41, 8)),
	3517 => std_logic_vector(to_unsigned(41, 8)),
	3518 => std_logic_vector(to_unsigned(42, 8)),
	3519 => std_logic_vector(to_unsigned(41, 8)),
	3520 => std_logic_vector(to_unsigned(42, 8)),
	3521 => std_logic_vector(to_unsigned(41, 8)),
	3522 => std_logic_vector(to_unsigned(41, 8)),
	3523 => std_logic_vector(to_unsigned(42, 8)),
	3524 => std_logic_vector(to_unsigned(41, 8)),
	3525 => std_logic_vector(to_unsigned(42, 8)),
	3526 => std_logic_vector(to_unsigned(42, 8)),
	3527 => std_logic_vector(to_unsigned(42, 8)),
	3528 => std_logic_vector(to_unsigned(42, 8)),
	3529 => std_logic_vector(to_unsigned(42, 8)),
	3530 => std_logic_vector(to_unsigned(41, 8)),
	3531 => std_logic_vector(to_unsigned(42, 8)),
	3532 => std_logic_vector(to_unsigned(41, 8)),
	3533 => std_logic_vector(to_unsigned(42, 8)),
	3534 => std_logic_vector(to_unsigned(42, 8)),
	3535 => std_logic_vector(to_unsigned(41, 8)),
	3536 => std_logic_vector(to_unsigned(42, 8)),
	3537 => std_logic_vector(to_unsigned(42, 8)),
	3538 => std_logic_vector(to_unsigned(42, 8)),
	3539 => std_logic_vector(to_unsigned(41, 8)),
	3540 => std_logic_vector(to_unsigned(41, 8)),
	3541 => std_logic_vector(to_unsigned(41, 8)),
	3542 => std_logic_vector(to_unsigned(42, 8)),
	3543 => std_logic_vector(to_unsigned(42, 8)),
	3544 => std_logic_vector(to_unsigned(42, 8)),
	3545 => std_logic_vector(to_unsigned(42, 8)),
	3546 => std_logic_vector(to_unsigned(41, 8)),
	3547 => std_logic_vector(to_unsigned(41, 8)),
	3548 => std_logic_vector(to_unsigned(41, 8)),
	3549 => std_logic_vector(to_unsigned(42, 8)),
	3550 => std_logic_vector(to_unsigned(42, 8)),
	3551 => std_logic_vector(to_unsigned(41, 8)),
	3552 => std_logic_vector(to_unsigned(42, 8)),
	3553 => std_logic_vector(to_unsigned(41, 8)),
	3554 => std_logic_vector(to_unsigned(41, 8)),
	3555 => std_logic_vector(to_unsigned(42, 8)),
	3556 => std_logic_vector(to_unsigned(42, 8)),
	3557 => std_logic_vector(to_unsigned(42, 8)),
	3558 => std_logic_vector(to_unsigned(42, 8)),
	3559 => std_logic_vector(to_unsigned(42, 8)),
	3560 => std_logic_vector(to_unsigned(42, 8)),
	3561 => std_logic_vector(to_unsigned(41, 8)),
	3562 => std_logic_vector(to_unsigned(42, 8)),
	3563 => std_logic_vector(to_unsigned(41, 8)),
	3564 => std_logic_vector(to_unsigned(41, 8)),
	3565 => std_logic_vector(to_unsigned(41, 8)),
	3566 => std_logic_vector(to_unsigned(42, 8)),
	3567 => std_logic_vector(to_unsigned(41, 8)),
	3568 => std_logic_vector(to_unsigned(42, 8)),
	3569 => std_logic_vector(to_unsigned(42, 8)),
	3570 => std_logic_vector(to_unsigned(42, 8)),
	3571 => std_logic_vector(to_unsigned(42, 8)),
	3572 => std_logic_vector(to_unsigned(42, 8)),
	3573 => std_logic_vector(to_unsigned(41, 8)),
	3574 => std_logic_vector(to_unsigned(41, 8)),
	3575 => std_logic_vector(to_unsigned(41, 8)),
	3576 => std_logic_vector(to_unsigned(42, 8)),
	3577 => std_logic_vector(to_unsigned(42, 8)),
	3578 => std_logic_vector(to_unsigned(41, 8)),
	3579 => std_logic_vector(to_unsigned(42, 8)),
	3580 => std_logic_vector(to_unsigned(42, 8)),
	3581 => std_logic_vector(to_unsigned(42, 8)),
	3582 => std_logic_vector(to_unsigned(42, 8)),
	3583 => std_logic_vector(to_unsigned(42, 8)),
	3584 => std_logic_vector(to_unsigned(41, 8)),
	3585 => std_logic_vector(to_unsigned(42, 8)),
	3586 => std_logic_vector(to_unsigned(41, 8)),
	3587 => std_logic_vector(to_unsigned(41, 8)),
	3588 => std_logic_vector(to_unsigned(41, 8)),
	3589 => std_logic_vector(to_unsigned(42, 8)),
	3590 => std_logic_vector(to_unsigned(41, 8)),
	3591 => std_logic_vector(to_unsigned(42, 8)),
	3592 => std_logic_vector(to_unsigned(42, 8)),
	3593 => std_logic_vector(to_unsigned(42, 8)),
	3594 => std_logic_vector(to_unsigned(41, 8)),
	3595 => std_logic_vector(to_unsigned(41, 8)),
	3596 => std_logic_vector(to_unsigned(41, 8)),
	3597 => std_logic_vector(to_unsigned(41, 8)),
	3598 => std_logic_vector(to_unsigned(42, 8)),
	3599 => std_logic_vector(to_unsigned(41, 8)),
	3600 => std_logic_vector(to_unsigned(41, 8)),
	3601 => std_logic_vector(to_unsigned(41, 8)),
	3602 => std_logic_vector(to_unsigned(41, 8)),
	3603 => std_logic_vector(to_unsigned(41, 8)),
	3604 => std_logic_vector(to_unsigned(42, 8)),
	3605 => std_logic_vector(to_unsigned(41, 8)),
	3606 => std_logic_vector(to_unsigned(42, 8)),
	3607 => std_logic_vector(to_unsigned(41, 8)),
	3608 => std_logic_vector(to_unsigned(41, 8)),
	3609 => std_logic_vector(to_unsigned(41, 8)),
	3610 => std_logic_vector(to_unsigned(42, 8)),
	3611 => std_logic_vector(to_unsigned(42, 8)),
	3612 => std_logic_vector(to_unsigned(42, 8)),
	3613 => std_logic_vector(to_unsigned(42, 8)),
	3614 => std_logic_vector(to_unsigned(41, 8)),
	3615 => std_logic_vector(to_unsigned(41, 8)),
	3616 => std_logic_vector(to_unsigned(42, 8)),
	3617 => std_logic_vector(to_unsigned(42, 8)),
	3618 => std_logic_vector(to_unsigned(42, 8)),
	3619 => std_logic_vector(to_unsigned(42, 8)),
	3620 => std_logic_vector(to_unsigned(41, 8)),
	3621 => std_logic_vector(to_unsigned(41, 8)),
	3622 => std_logic_vector(to_unsigned(41, 8)),
	3623 => std_logic_vector(to_unsigned(42, 8)),
	3624 => std_logic_vector(to_unsigned(42, 8)),
	3625 => std_logic_vector(to_unsigned(41, 8)),
	3626 => std_logic_vector(to_unsigned(42, 8)),
	3627 => std_logic_vector(to_unsigned(42, 8)),
	3628 => std_logic_vector(to_unsigned(41, 8)),
	3629 => std_logic_vector(to_unsigned(41, 8)),
	3630 => std_logic_vector(to_unsigned(41, 8)),
	3631 => std_logic_vector(to_unsigned(41, 8)),
	3632 => std_logic_vector(to_unsigned(42, 8)),
	3633 => std_logic_vector(to_unsigned(41, 8)),
	3634 => std_logic_vector(to_unsigned(41, 8)),
	3635 => std_logic_vector(to_unsigned(41, 8)),
	3636 => std_logic_vector(to_unsigned(42, 8)),
	3637 => std_logic_vector(to_unsigned(42, 8)),
	3638 => std_logic_vector(to_unsigned(42, 8)),
	3639 => std_logic_vector(to_unsigned(42, 8)),
	3640 => std_logic_vector(to_unsigned(41, 8)),
	3641 => std_logic_vector(to_unsigned(42, 8)),
	3642 => std_logic_vector(to_unsigned(41, 8)),
	3643 => std_logic_vector(to_unsigned(42, 8)),
	3644 => std_logic_vector(to_unsigned(41, 8)),
	3645 => std_logic_vector(to_unsigned(42, 8)),
	3646 => std_logic_vector(to_unsigned(42, 8)),
	3647 => std_logic_vector(to_unsigned(41, 8)),
	3648 => std_logic_vector(to_unsigned(41, 8)),
	3649 => std_logic_vector(to_unsigned(41, 8)),
	3650 => std_logic_vector(to_unsigned(41, 8)),
	3651 => std_logic_vector(to_unsigned(41, 8)),
	3652 => std_logic_vector(to_unsigned(41, 8)),
	3653 => std_logic_vector(to_unsigned(41, 8)),
	3654 => std_logic_vector(to_unsigned(42, 8)),
	3655 => std_logic_vector(to_unsigned(42, 8)),
	3656 => std_logic_vector(to_unsigned(42, 8)),
	3657 => std_logic_vector(to_unsigned(42, 8)),
	3658 => std_logic_vector(to_unsigned(41, 8)),
	3659 => std_logic_vector(to_unsigned(41, 8)),
	3660 => std_logic_vector(to_unsigned(41, 8)),
	3661 => std_logic_vector(to_unsigned(41, 8)),
	3662 => std_logic_vector(to_unsigned(41, 8)),
	3663 => std_logic_vector(to_unsigned(41, 8)),
	3664 => std_logic_vector(to_unsigned(41, 8)),
	3665 => std_logic_vector(to_unsigned(42, 8)),
	3666 => std_logic_vector(to_unsigned(42, 8)),
	3667 => std_logic_vector(to_unsigned(41, 8)),
	3668 => std_logic_vector(to_unsigned(41, 8)),
	3669 => std_logic_vector(to_unsigned(41, 8)),
	3670 => std_logic_vector(to_unsigned(42, 8)),
	3671 => std_logic_vector(to_unsigned(42, 8)),
	3672 => std_logic_vector(to_unsigned(41, 8)),
	3673 => std_logic_vector(to_unsigned(41, 8)),
	3674 => std_logic_vector(to_unsigned(41, 8)),
	3675 => std_logic_vector(to_unsigned(42, 8)),
	3676 => std_logic_vector(to_unsigned(41, 8)),
	3677 => std_logic_vector(to_unsigned(41, 8)),
	3678 => std_logic_vector(to_unsigned(41, 8)),
	3679 => std_logic_vector(to_unsigned(42, 8)),
	3680 => std_logic_vector(to_unsigned(42, 8)),
	3681 => std_logic_vector(to_unsigned(42, 8)),
	3682 => std_logic_vector(to_unsigned(41, 8)),
	3683 => std_logic_vector(to_unsigned(42, 8)),
	3684 => std_logic_vector(to_unsigned(41, 8)),
	3685 => std_logic_vector(to_unsigned(41, 8)),
	3686 => std_logic_vector(to_unsigned(42, 8)),
	3687 => std_logic_vector(to_unsigned(42, 8)),
	3688 => std_logic_vector(to_unsigned(42, 8)),
	3689 => std_logic_vector(to_unsigned(41, 8)),
	3690 => std_logic_vector(to_unsigned(42, 8)),
	3691 => std_logic_vector(to_unsigned(41, 8)),
	3692 => std_logic_vector(to_unsigned(41, 8)),
	3693 => std_logic_vector(to_unsigned(42, 8)),
	3694 => std_logic_vector(to_unsigned(41, 8)),
	3695 => std_logic_vector(to_unsigned(42, 8)),
	3696 => std_logic_vector(to_unsigned(42, 8)),
	3697 => std_logic_vector(to_unsigned(42, 8)),
	3698 => std_logic_vector(to_unsigned(42, 8)),
	3699 => std_logic_vector(to_unsigned(42, 8)),
	3700 => std_logic_vector(to_unsigned(42, 8)),
	3701 => std_logic_vector(to_unsigned(41, 8)),
	3702 => std_logic_vector(to_unsigned(41, 8)),
	3703 => std_logic_vector(to_unsigned(42, 8)),
	3704 => std_logic_vector(to_unsigned(41, 8)),
	3705 => std_logic_vector(to_unsigned(41, 8)),
	3706 => std_logic_vector(to_unsigned(41, 8)),
	3707 => std_logic_vector(to_unsigned(42, 8)),
	3708 => std_logic_vector(to_unsigned(41, 8)),
	3709 => std_logic_vector(to_unsigned(42, 8)),
	3710 => std_logic_vector(to_unsigned(42, 8)),
	3711 => std_logic_vector(to_unsigned(41, 8)),
	3712 => std_logic_vector(to_unsigned(42, 8)),
	3713 => std_logic_vector(to_unsigned(42, 8)),
	3714 => std_logic_vector(to_unsigned(42, 8)),
	3715 => std_logic_vector(to_unsigned(41, 8)),
	3716 => std_logic_vector(to_unsigned(42, 8)),
	3717 => std_logic_vector(to_unsigned(42, 8)),
	3718 => std_logic_vector(to_unsigned(42, 8)),
	3719 => std_logic_vector(to_unsigned(42, 8)),
	3720 => std_logic_vector(to_unsigned(42, 8)),
	3721 => std_logic_vector(to_unsigned(42, 8)),
	3722 => std_logic_vector(to_unsigned(42, 8)),
	3723 => std_logic_vector(to_unsigned(41, 8)),
	3724 => std_logic_vector(to_unsigned(41, 8)),
	3725 => std_logic_vector(to_unsigned(42, 8)),
	3726 => std_logic_vector(to_unsigned(42, 8)),
	3727 => std_logic_vector(to_unsigned(41, 8)),
	3728 => std_logic_vector(to_unsigned(42, 8)),
	3729 => std_logic_vector(to_unsigned(42, 8)),
	3730 => std_logic_vector(to_unsigned(42, 8)),
	3731 => std_logic_vector(to_unsigned(42, 8)),
	3732 => std_logic_vector(to_unsigned(42, 8)),
	3733 => std_logic_vector(to_unsigned(41, 8)),
	3734 => std_logic_vector(to_unsigned(41, 8)),
	3735 => std_logic_vector(to_unsigned(41, 8)),
	3736 => std_logic_vector(to_unsigned(41, 8)),
	3737 => std_logic_vector(to_unsigned(42, 8)),
	3738 => std_logic_vector(to_unsigned(42, 8)),
	3739 => std_logic_vector(to_unsigned(42, 8)),
	3740 => std_logic_vector(to_unsigned(41, 8)),
	3741 => std_logic_vector(to_unsigned(41, 8)),
	3742 => std_logic_vector(to_unsigned(41, 8)),
	3743 => std_logic_vector(to_unsigned(42, 8)),
	3744 => std_logic_vector(to_unsigned(42, 8)),
	3745 => std_logic_vector(to_unsigned(42, 8)),
	3746 => std_logic_vector(to_unsigned(42, 8)),
	3747 => std_logic_vector(to_unsigned(42, 8)),
	3748 => std_logic_vector(to_unsigned(41, 8)),
	3749 => std_logic_vector(to_unsigned(42, 8)),
	3750 => std_logic_vector(to_unsigned(42, 8)),
	3751 => std_logic_vector(to_unsigned(42, 8)),
	3752 => std_logic_vector(to_unsigned(41, 8)),
	3753 => std_logic_vector(to_unsigned(42, 8)),
	3754 => std_logic_vector(to_unsigned(41, 8)),
	3755 => std_logic_vector(to_unsigned(42, 8)),
	3756 => std_logic_vector(to_unsigned(41, 8)),
	3757 => std_logic_vector(to_unsigned(42, 8)),
	3758 => std_logic_vector(to_unsigned(41, 8)),
	3759 => std_logic_vector(to_unsigned(41, 8)),
	3760 => std_logic_vector(to_unsigned(41, 8)),
	3761 => std_logic_vector(to_unsigned(42, 8)),
	3762 => std_logic_vector(to_unsigned(42, 8)),
	3763 => std_logic_vector(to_unsigned(41, 8)),
	3764 => std_logic_vector(to_unsigned(42, 8)),
	3765 => std_logic_vector(to_unsigned(41, 8)),
	3766 => std_logic_vector(to_unsigned(42, 8)),
	3767 => std_logic_vector(to_unsigned(41, 8)),
	3768 => std_logic_vector(to_unsigned(41, 8)),
	3769 => std_logic_vector(to_unsigned(42, 8)),
	3770 => std_logic_vector(to_unsigned(42, 8)),
	3771 => std_logic_vector(to_unsigned(41, 8)),
	3772 => std_logic_vector(to_unsigned(41, 8)),
	3773 => std_logic_vector(to_unsigned(42, 8)),
	3774 => std_logic_vector(to_unsigned(42, 8)),
	3775 => std_logic_vector(to_unsigned(42, 8)),
	3776 => std_logic_vector(to_unsigned(41, 8)),
	3777 => std_logic_vector(to_unsigned(42, 8)),
	3778 => std_logic_vector(to_unsigned(42, 8)),
	3779 => std_logic_vector(to_unsigned(41, 8)),
	3780 => std_logic_vector(to_unsigned(42, 8)),
	3781 => std_logic_vector(to_unsigned(42, 8)),
	3782 => std_logic_vector(to_unsigned(41, 8)),
	3783 => std_logic_vector(to_unsigned(42, 8)),
	3784 => std_logic_vector(to_unsigned(42, 8)),
	3785 => std_logic_vector(to_unsigned(41, 8)),
	3786 => std_logic_vector(to_unsigned(42, 8)),
	3787 => std_logic_vector(to_unsigned(41, 8)),
	3788 => std_logic_vector(to_unsigned(42, 8)),
	3789 => std_logic_vector(to_unsigned(41, 8)),
	3790 => std_logic_vector(to_unsigned(42, 8)),
	3791 => std_logic_vector(to_unsigned(42, 8)),
	3792 => std_logic_vector(to_unsigned(42, 8)),
	3793 => std_logic_vector(to_unsigned(41, 8)),
	3794 => std_logic_vector(to_unsigned(41, 8)),
	3795 => std_logic_vector(to_unsigned(42, 8)),
	3796 => std_logic_vector(to_unsigned(42, 8)),
	3797 => std_logic_vector(to_unsigned(42, 8)),
	3798 => std_logic_vector(to_unsigned(41, 8)),
	3799 => std_logic_vector(to_unsigned(42, 8)),
	3800 => std_logic_vector(to_unsigned(41, 8)),
	3801 => std_logic_vector(to_unsigned(41, 8)),
	3802 => std_logic_vector(to_unsigned(41, 8)),
	3803 => std_logic_vector(to_unsigned(42, 8)),
	3804 => std_logic_vector(to_unsigned(42, 8)),
	3805 => std_logic_vector(to_unsigned(42, 8)),
	3806 => std_logic_vector(to_unsigned(41, 8)),
	3807 => std_logic_vector(to_unsigned(42, 8)),
	3808 => std_logic_vector(to_unsigned(42, 8)),
	3809 => std_logic_vector(to_unsigned(41, 8)),
	3810 => std_logic_vector(to_unsigned(42, 8)),
	3811 => std_logic_vector(to_unsigned(41, 8)),
	3812 => std_logic_vector(to_unsigned(42, 8)),
	3813 => std_logic_vector(to_unsigned(41, 8)),
	3814 => std_logic_vector(to_unsigned(41, 8)),
	3815 => std_logic_vector(to_unsigned(42, 8)),
	3816 => std_logic_vector(to_unsigned(41, 8)),
	3817 => std_logic_vector(to_unsigned(41, 8)),
	3818 => std_logic_vector(to_unsigned(42, 8)),
	3819 => std_logic_vector(to_unsigned(42, 8)),
	3820 => std_logic_vector(to_unsigned(41, 8)),
	3821 => std_logic_vector(to_unsigned(41, 8)),
	3822 => std_logic_vector(to_unsigned(42, 8)),
	3823 => std_logic_vector(to_unsigned(42, 8)),
	3824 => std_logic_vector(to_unsigned(41, 8)),
	3825 => std_logic_vector(to_unsigned(41, 8)),
	3826 => std_logic_vector(to_unsigned(42, 8)),
	3827 => std_logic_vector(to_unsigned(42, 8)),
	3828 => std_logic_vector(to_unsigned(41, 8)),
	3829 => std_logic_vector(to_unsigned(41, 8)),
	3830 => std_logic_vector(to_unsigned(42, 8)),
	3831 => std_logic_vector(to_unsigned(42, 8)),
	3832 => std_logic_vector(to_unsigned(42, 8)),
	3833 => std_logic_vector(to_unsigned(41, 8)),
	3834 => std_logic_vector(to_unsigned(42, 8)),
	3835 => std_logic_vector(to_unsigned(42, 8)),
	3836 => std_logic_vector(to_unsigned(41, 8)),
	3837 => std_logic_vector(to_unsigned(41, 8)),
	3838 => std_logic_vector(to_unsigned(41, 8)),
	3839 => std_logic_vector(to_unsigned(41, 8)),
	3840 => std_logic_vector(to_unsigned(42, 8)),
	3841 => std_logic_vector(to_unsigned(41, 8)),
	3842 => std_logic_vector(to_unsigned(41, 8)),
	3843 => std_logic_vector(to_unsigned(42, 8)),
	3844 => std_logic_vector(to_unsigned(41, 8)),
	3845 => std_logic_vector(to_unsigned(42, 8)),
	3846 => std_logic_vector(to_unsigned(42, 8)),
	3847 => std_logic_vector(to_unsigned(42, 8)),
	3848 => std_logic_vector(to_unsigned(42, 8)),
	3849 => std_logic_vector(to_unsigned(42, 8)),
	3850 => std_logic_vector(to_unsigned(42, 8)),
	3851 => std_logic_vector(to_unsigned(42, 8)),
	3852 => std_logic_vector(to_unsigned(41, 8)),
	3853 => std_logic_vector(to_unsigned(42, 8)),
	3854 => std_logic_vector(to_unsigned(42, 8)),
	3855 => std_logic_vector(to_unsigned(42, 8)),
	3856 => std_logic_vector(to_unsigned(41, 8)),
	3857 => std_logic_vector(to_unsigned(42, 8)),
	3858 => std_logic_vector(to_unsigned(42, 8)),
	3859 => std_logic_vector(to_unsigned(41, 8)),
	3860 => std_logic_vector(to_unsigned(41, 8)),
	3861 => std_logic_vector(to_unsigned(42, 8)),
	3862 => std_logic_vector(to_unsigned(42, 8)),
	3863 => std_logic_vector(to_unsigned(42, 8)),
	3864 => std_logic_vector(to_unsigned(42, 8)),
	3865 => std_logic_vector(to_unsigned(42, 8)),
	3866 => std_logic_vector(to_unsigned(42, 8)),
	3867 => std_logic_vector(to_unsigned(41, 8)),
	3868 => std_logic_vector(to_unsigned(42, 8)),
	3869 => std_logic_vector(to_unsigned(42, 8)),
	3870 => std_logic_vector(to_unsigned(42, 8)),
	3871 => std_logic_vector(to_unsigned(42, 8)),
	3872 => std_logic_vector(to_unsigned(41, 8)),
	3873 => std_logic_vector(to_unsigned(41, 8)),
	3874 => std_logic_vector(to_unsigned(42, 8)),
	3875 => std_logic_vector(to_unsigned(42, 8)),
	3876 => std_logic_vector(to_unsigned(42, 8)),
	3877 => std_logic_vector(to_unsigned(41, 8)),
	3878 => std_logic_vector(to_unsigned(41, 8)),
	3879 => std_logic_vector(to_unsigned(42, 8)),
	3880 => std_logic_vector(to_unsigned(42, 8)),
	3881 => std_logic_vector(to_unsigned(42, 8)),
	3882 => std_logic_vector(to_unsigned(42, 8)),
	3883 => std_logic_vector(to_unsigned(42, 8)),
	3884 => std_logic_vector(to_unsigned(42, 8)),
	3885 => std_logic_vector(to_unsigned(41, 8)),
	3886 => std_logic_vector(to_unsigned(42, 8)),
	3887 => std_logic_vector(to_unsigned(41, 8)),
	3888 => std_logic_vector(to_unsigned(42, 8)),
	3889 => std_logic_vector(to_unsigned(41, 8)),
	3890 => std_logic_vector(to_unsigned(41, 8)),
	3891 => std_logic_vector(to_unsigned(41, 8)),
	3892 => std_logic_vector(to_unsigned(41, 8)),
	3893 => std_logic_vector(to_unsigned(41, 8)),
	3894 => std_logic_vector(to_unsigned(41, 8)),
	3895 => std_logic_vector(to_unsigned(42, 8)),
	3896 => std_logic_vector(to_unsigned(41, 8)),
	3897 => std_logic_vector(to_unsigned(41, 8)),
	3898 => std_logic_vector(to_unsigned(41, 8)),
	3899 => std_logic_vector(to_unsigned(41, 8)),
	3900 => std_logic_vector(to_unsigned(41, 8)),
	3901 => std_logic_vector(to_unsigned(41, 8)),
	3902 => std_logic_vector(to_unsigned(41, 8)),
	3903 => std_logic_vector(to_unsigned(42, 8)),
	3904 => std_logic_vector(to_unsigned(41, 8)),
	3905 => std_logic_vector(to_unsigned(42, 8)),
	3906 => std_logic_vector(to_unsigned(42, 8)),
	3907 => std_logic_vector(to_unsigned(42, 8)),
	3908 => std_logic_vector(to_unsigned(41, 8)),
	3909 => std_logic_vector(to_unsigned(41, 8)),
	3910 => std_logic_vector(to_unsigned(42, 8)),
	3911 => std_logic_vector(to_unsigned(42, 8)),
	3912 => std_logic_vector(to_unsigned(41, 8)),
	3913 => std_logic_vector(to_unsigned(42, 8)),
	3914 => std_logic_vector(to_unsigned(42, 8)),
	3915 => std_logic_vector(to_unsigned(41, 8)),
	3916 => std_logic_vector(to_unsigned(41, 8)),
	3917 => std_logic_vector(to_unsigned(42, 8)),
	3918 => std_logic_vector(to_unsigned(42, 8)),
	3919 => std_logic_vector(to_unsigned(42, 8)),
	3920 => std_logic_vector(to_unsigned(42, 8)),
	3921 => std_logic_vector(to_unsigned(41, 8)),
	3922 => std_logic_vector(to_unsigned(41, 8)),
	3923 => std_logic_vector(to_unsigned(42, 8)),
	3924 => std_logic_vector(to_unsigned(42, 8)),
	3925 => std_logic_vector(to_unsigned(42, 8)),
	3926 => std_logic_vector(to_unsigned(41, 8)),
	3927 => std_logic_vector(to_unsigned(41, 8)),
	3928 => std_logic_vector(to_unsigned(42, 8)),
	3929 => std_logic_vector(to_unsigned(42, 8)),
	3930 => std_logic_vector(to_unsigned(41, 8)),
	3931 => std_logic_vector(to_unsigned(42, 8)),
	3932 => std_logic_vector(to_unsigned(42, 8)),
	3933 => std_logic_vector(to_unsigned(42, 8)),
	3934 => std_logic_vector(to_unsigned(41, 8)),
	3935 => std_logic_vector(to_unsigned(42, 8)),
	3936 => std_logic_vector(to_unsigned(41, 8)),
	3937 => std_logic_vector(to_unsigned(41, 8)),
	3938 => std_logic_vector(to_unsigned(41, 8)),
	3939 => std_logic_vector(to_unsigned(41, 8)),
	3940 => std_logic_vector(to_unsigned(41, 8)),
	3941 => std_logic_vector(to_unsigned(42, 8)),
	3942 => std_logic_vector(to_unsigned(42, 8)),
	3943 => std_logic_vector(to_unsigned(41, 8)),
	3944 => std_logic_vector(to_unsigned(41, 8)),
	3945 => std_logic_vector(to_unsigned(42, 8)),
	3946 => std_logic_vector(to_unsigned(41, 8)),
	3947 => std_logic_vector(to_unsigned(42, 8)),
	3948 => std_logic_vector(to_unsigned(41, 8)),
	3949 => std_logic_vector(to_unsigned(42, 8)),
	3950 => std_logic_vector(to_unsigned(42, 8)),
	3951 => std_logic_vector(to_unsigned(41, 8)),
	3952 => std_logic_vector(to_unsigned(42, 8)),
	3953 => std_logic_vector(to_unsigned(41, 8)),
	3954 => std_logic_vector(to_unsigned(42, 8)),
	3955 => std_logic_vector(to_unsigned(41, 8)),
	3956 => std_logic_vector(to_unsigned(42, 8)),
	3957 => std_logic_vector(to_unsigned(41, 8)),
	3958 => std_logic_vector(to_unsigned(42, 8)),
	3959 => std_logic_vector(to_unsigned(42, 8)),
	3960 => std_logic_vector(to_unsigned(42, 8)),
	3961 => std_logic_vector(to_unsigned(41, 8)),
	3962 => std_logic_vector(to_unsigned(41, 8)),
	3963 => std_logic_vector(to_unsigned(41, 8)),
	3964 => std_logic_vector(to_unsigned(42, 8)),
	3965 => std_logic_vector(to_unsigned(42, 8)),
	3966 => std_logic_vector(to_unsigned(41, 8)),
	3967 => std_logic_vector(to_unsigned(41, 8)),
	3968 => std_logic_vector(to_unsigned(41, 8)),
	3969 => std_logic_vector(to_unsigned(41, 8)),
	3970 => std_logic_vector(to_unsigned(42, 8)),
	3971 => std_logic_vector(to_unsigned(41, 8)),
	3972 => std_logic_vector(to_unsigned(41, 8)),
	3973 => std_logic_vector(to_unsigned(41, 8)),
	3974 => std_logic_vector(to_unsigned(41, 8)),
	3975 => std_logic_vector(to_unsigned(41, 8)),
	3976 => std_logic_vector(to_unsigned(41, 8)),
	3977 => std_logic_vector(to_unsigned(42, 8)),
	3978 => std_logic_vector(to_unsigned(41, 8)),
	3979 => std_logic_vector(to_unsigned(42, 8)),
	3980 => std_logic_vector(to_unsigned(41, 8)),
	3981 => std_logic_vector(to_unsigned(42, 8)),
	3982 => std_logic_vector(to_unsigned(42, 8)),
	3983 => std_logic_vector(to_unsigned(41, 8)),
	3984 => std_logic_vector(to_unsigned(42, 8)),
	3985 => std_logic_vector(to_unsigned(41, 8)),
	3986 => std_logic_vector(to_unsigned(42, 8)),
	3987 => std_logic_vector(to_unsigned(41, 8)),
	3988 => std_logic_vector(to_unsigned(41, 8)),
	3989 => std_logic_vector(to_unsigned(41, 8)),
	3990 => std_logic_vector(to_unsigned(42, 8)),
	3991 => std_logic_vector(to_unsigned(41, 8)),
	3992 => std_logic_vector(to_unsigned(42, 8)),
	3993 => std_logic_vector(to_unsigned(41, 8)),
	3994 => std_logic_vector(to_unsigned(41, 8)),
	3995 => std_logic_vector(to_unsigned(41, 8)),
	3996 => std_logic_vector(to_unsigned(41, 8)),
	3997 => std_logic_vector(to_unsigned(42, 8)),
	3998 => std_logic_vector(to_unsigned(42, 8)),
	3999 => std_logic_vector(to_unsigned(42, 8)),
	4000 => std_logic_vector(to_unsigned(42, 8)),
	4001 => std_logic_vector(to_unsigned(42, 8)),
	4002 => std_logic_vector(to_unsigned(41, 8)),
	4003 => std_logic_vector(to_unsigned(42, 8)),
	4004 => std_logic_vector(to_unsigned(41, 8)),
	4005 => std_logic_vector(to_unsigned(42, 8)),
	4006 => std_logic_vector(to_unsigned(41, 8)),
	4007 => std_logic_vector(to_unsigned(42, 8)),
	4008 => std_logic_vector(to_unsigned(41, 8)),
	4009 => std_logic_vector(to_unsigned(42, 8)),
	4010 => std_logic_vector(to_unsigned(41, 8)),
	4011 => std_logic_vector(to_unsigned(41, 8)),
	4012 => std_logic_vector(to_unsigned(42, 8)),
	4013 => std_logic_vector(to_unsigned(41, 8)),
	4014 => std_logic_vector(to_unsigned(41, 8)),
	4015 => std_logic_vector(to_unsigned(42, 8)),
	4016 => std_logic_vector(to_unsigned(42, 8)),
	4017 => std_logic_vector(to_unsigned(42, 8)),
	4018 => std_logic_vector(to_unsigned(41, 8)),
	4019 => std_logic_vector(to_unsigned(41, 8)),
	4020 => std_logic_vector(to_unsigned(41, 8)),
	4021 => std_logic_vector(to_unsigned(41, 8)),
	4022 => std_logic_vector(to_unsigned(42, 8)),
	4023 => std_logic_vector(to_unsigned(41, 8)),
	4024 => std_logic_vector(to_unsigned(42, 8)),
	4025 => std_logic_vector(to_unsigned(41, 8)),
	4026 => std_logic_vector(to_unsigned(41, 8)),
	4027 => std_logic_vector(to_unsigned(41, 8)),
	4028 => std_logic_vector(to_unsigned(41, 8)),
	4029 => std_logic_vector(to_unsigned(42, 8)),
	4030 => std_logic_vector(to_unsigned(42, 8)),
	4031 => std_logic_vector(to_unsigned(41, 8)),
	4032 => std_logic_vector(to_unsigned(41, 8)),
	4033 => std_logic_vector(to_unsigned(42, 8)),
	4034 => std_logic_vector(to_unsigned(41, 8)),
	4035 => std_logic_vector(to_unsigned(42, 8)),
	4036 => std_logic_vector(to_unsigned(41, 8)),
	4037 => std_logic_vector(to_unsigned(42, 8)),
	4038 => std_logic_vector(to_unsigned(42, 8)),
	4039 => std_logic_vector(to_unsigned(41, 8)),
	4040 => std_logic_vector(to_unsigned(42, 8)),
	4041 => std_logic_vector(to_unsigned(42, 8)),
	4042 => std_logic_vector(to_unsigned(42, 8)),
	4043 => std_logic_vector(to_unsigned(41, 8)),
	4044 => std_logic_vector(to_unsigned(41, 8)),
	4045 => std_logic_vector(to_unsigned(42, 8)),
	4046 => std_logic_vector(to_unsigned(42, 8)),
	4047 => std_logic_vector(to_unsigned(42, 8)),
	4048 => std_logic_vector(to_unsigned(41, 8)),
	4049 => std_logic_vector(to_unsigned(42, 8)),
	4050 => std_logic_vector(to_unsigned(42, 8)),
	4051 => std_logic_vector(to_unsigned(41, 8)),
	4052 => std_logic_vector(to_unsigned(42, 8)),
	4053 => std_logic_vector(to_unsigned(41, 8)),
	4054 => std_logic_vector(to_unsigned(42, 8)),
	4055 => std_logic_vector(to_unsigned(41, 8)),
	4056 => std_logic_vector(to_unsigned(42, 8)),
	4057 => std_logic_vector(to_unsigned(42, 8)),
	4058 => std_logic_vector(to_unsigned(41, 8)),
	4059 => std_logic_vector(to_unsigned(42, 8)),
	4060 => std_logic_vector(to_unsigned(42, 8)),
	4061 => std_logic_vector(to_unsigned(42, 8)),
	4062 => std_logic_vector(to_unsigned(42, 8)),
	4063 => std_logic_vector(to_unsigned(41, 8)),
	4064 => std_logic_vector(to_unsigned(41, 8)),
	4065 => std_logic_vector(to_unsigned(41, 8)),
	4066 => std_logic_vector(to_unsigned(42, 8)),
	4067 => std_logic_vector(to_unsigned(41, 8)),
	4068 => std_logic_vector(to_unsigned(42, 8)),
	4069 => std_logic_vector(to_unsigned(42, 8)),
	4070 => std_logic_vector(to_unsigned(42, 8)),
	4071 => std_logic_vector(to_unsigned(42, 8)),
	4072 => std_logic_vector(to_unsigned(41, 8)),
	4073 => std_logic_vector(to_unsigned(41, 8)),
	4074 => std_logic_vector(to_unsigned(41, 8)),
	4075 => std_logic_vector(to_unsigned(41, 8)),
	4076 => std_logic_vector(to_unsigned(41, 8)),
	4077 => std_logic_vector(to_unsigned(41, 8)),
	4078 => std_logic_vector(to_unsigned(41, 8)),
	4079 => std_logic_vector(to_unsigned(41, 8)),
	4080 => std_logic_vector(to_unsigned(42, 8)),
	4081 => std_logic_vector(to_unsigned(42, 8)),
	4082 => std_logic_vector(to_unsigned(42, 8)),
	4083 => std_logic_vector(to_unsigned(42, 8)),
	4084 => std_logic_vector(to_unsigned(42, 8)),
	4085 => std_logic_vector(to_unsigned(41, 8)),
	4086 => std_logic_vector(to_unsigned(42, 8)),
	4087 => std_logic_vector(to_unsigned(41, 8)),
	4088 => std_logic_vector(to_unsigned(41, 8)),
	4089 => std_logic_vector(to_unsigned(41, 8)),
	4090 => std_logic_vector(to_unsigned(42, 8)),
	4091 => std_logic_vector(to_unsigned(41, 8)),
	4092 => std_logic_vector(to_unsigned(41, 8)),
	4093 => std_logic_vector(to_unsigned(41, 8)),
	4094 => std_logic_vector(to_unsigned(42, 8)),
	4095 => std_logic_vector(to_unsigned(41, 8)),
	4096 => std_logic_vector(to_unsigned(41, 8)),
	4097 => std_logic_vector(to_unsigned(42, 8)),
	4098 => std_logic_vector(to_unsigned(41, 8)),
	4099 => std_logic_vector(to_unsigned(41, 8)),
	4100 => std_logic_vector(to_unsigned(41, 8)),
	4101 => std_logic_vector(to_unsigned(42, 8)),
	4102 => std_logic_vector(to_unsigned(41, 8)),
	4103 => std_logic_vector(to_unsigned(42, 8)),
	4104 => std_logic_vector(to_unsigned(42, 8)),
	4105 => std_logic_vector(to_unsigned(41, 8)),
	4106 => std_logic_vector(to_unsigned(41, 8)),
	4107 => std_logic_vector(to_unsigned(42, 8)),
	4108 => std_logic_vector(to_unsigned(41, 8)),
	4109 => std_logic_vector(to_unsigned(41, 8)),
	4110 => std_logic_vector(to_unsigned(41, 8)),
	4111 => std_logic_vector(to_unsigned(42, 8)),
	4112 => std_logic_vector(to_unsigned(42, 8)),
	4113 => std_logic_vector(to_unsigned(42, 8)),
	4114 => std_logic_vector(to_unsigned(41, 8)),
	4115 => std_logic_vector(to_unsigned(41, 8)),
	4116 => std_logic_vector(to_unsigned(42, 8)),
	4117 => std_logic_vector(to_unsigned(42, 8)),
	4118 => std_logic_vector(to_unsigned(41, 8)),
	4119 => std_logic_vector(to_unsigned(42, 8)),
	4120 => std_logic_vector(to_unsigned(41, 8)),
	4121 => std_logic_vector(to_unsigned(42, 8)),
	4122 => std_logic_vector(to_unsigned(42, 8)),
	4123 => std_logic_vector(to_unsigned(42, 8)),
	4124 => std_logic_vector(to_unsigned(42, 8)),
	4125 => std_logic_vector(to_unsigned(41, 8)),
	4126 => std_logic_vector(to_unsigned(41, 8)),
	4127 => std_logic_vector(to_unsigned(42, 8)),
	4128 => std_logic_vector(to_unsigned(42, 8)),
	4129 => std_logic_vector(to_unsigned(42, 8)),
	4130 => std_logic_vector(to_unsigned(41, 8)),
	4131 => std_logic_vector(to_unsigned(42, 8)),
	4132 => std_logic_vector(to_unsigned(41, 8)),
	4133 => std_logic_vector(to_unsigned(42, 8)),
	4134 => std_logic_vector(to_unsigned(42, 8)),
	4135 => std_logic_vector(to_unsigned(41, 8)),
	4136 => std_logic_vector(to_unsigned(41, 8)),
	4137 => std_logic_vector(to_unsigned(41, 8)),
	4138 => std_logic_vector(to_unsigned(42, 8)),
	4139 => std_logic_vector(to_unsigned(41, 8)),
	4140 => std_logic_vector(to_unsigned(41, 8)),
	4141 => std_logic_vector(to_unsigned(42, 8)),
	4142 => std_logic_vector(to_unsigned(41, 8)),
	4143 => std_logic_vector(to_unsigned(42, 8)),
	4144 => std_logic_vector(to_unsigned(41, 8)),
	4145 => std_logic_vector(to_unsigned(42, 8)),
	4146 => std_logic_vector(to_unsigned(41, 8)),
	4147 => std_logic_vector(to_unsigned(42, 8)),
	4148 => std_logic_vector(to_unsigned(42, 8)),
	4149 => std_logic_vector(to_unsigned(41, 8)),
	4150 => std_logic_vector(to_unsigned(41, 8)),
	4151 => std_logic_vector(to_unsigned(42, 8)),
	4152 => std_logic_vector(to_unsigned(41, 8)),
	4153 => std_logic_vector(to_unsigned(41, 8)),
	4154 => std_logic_vector(to_unsigned(41, 8)),
	4155 => std_logic_vector(to_unsigned(42, 8)),
	4156 => std_logic_vector(to_unsigned(41, 8)),
	4157 => std_logic_vector(to_unsigned(41, 8)),
	4158 => std_logic_vector(to_unsigned(41, 8)),
	4159 => std_logic_vector(to_unsigned(42, 8)),
	4160 => std_logic_vector(to_unsigned(42, 8)),
	4161 => std_logic_vector(to_unsigned(42, 8)),
	4162 => std_logic_vector(to_unsigned(41, 8)),
	4163 => std_logic_vector(to_unsigned(41, 8)),
	4164 => std_logic_vector(to_unsigned(42, 8)),
	4165 => std_logic_vector(to_unsigned(41, 8)),
	4166 => std_logic_vector(to_unsigned(41, 8)),
	4167 => std_logic_vector(to_unsigned(42, 8)),
	4168 => std_logic_vector(to_unsigned(42, 8)),
	4169 => std_logic_vector(to_unsigned(41, 8)),
	4170 => std_logic_vector(to_unsigned(42, 8)),
	4171 => std_logic_vector(to_unsigned(42, 8)),
	4172 => std_logic_vector(to_unsigned(42, 8)),
	4173 => std_logic_vector(to_unsigned(41, 8)),
	4174 => std_logic_vector(to_unsigned(42, 8)),
	4175 => std_logic_vector(to_unsigned(42, 8)),
	4176 => std_logic_vector(to_unsigned(41, 8)),
	4177 => std_logic_vector(to_unsigned(42, 8)),
	4178 => std_logic_vector(to_unsigned(42, 8)),
	4179 => std_logic_vector(to_unsigned(41, 8)),
	4180 => std_logic_vector(to_unsigned(42, 8)),
	4181 => std_logic_vector(to_unsigned(41, 8)),
	4182 => std_logic_vector(to_unsigned(41, 8)),
	4183 => std_logic_vector(to_unsigned(41, 8)),
	4184 => std_logic_vector(to_unsigned(41, 8)),
	4185 => std_logic_vector(to_unsigned(42, 8)),
	4186 => std_logic_vector(to_unsigned(41, 8)),
	4187 => std_logic_vector(to_unsigned(41, 8)),
	4188 => std_logic_vector(to_unsigned(41, 8)),
	4189 => std_logic_vector(to_unsigned(41, 8)),
	4190 => std_logic_vector(to_unsigned(41, 8)),
	4191 => std_logic_vector(to_unsigned(41, 8)),
	4192 => std_logic_vector(to_unsigned(41, 8)),
	4193 => std_logic_vector(to_unsigned(42, 8)),
	4194 => std_logic_vector(to_unsigned(41, 8)),
	4195 => std_logic_vector(to_unsigned(42, 8)),
	4196 => std_logic_vector(to_unsigned(42, 8)),
	4197 => std_logic_vector(to_unsigned(42, 8)),
	4198 => std_logic_vector(to_unsigned(42, 8)),
	4199 => std_logic_vector(to_unsigned(42, 8)),
	4200 => std_logic_vector(to_unsigned(42, 8)),
	4201 => std_logic_vector(to_unsigned(41, 8)),
	4202 => std_logic_vector(to_unsigned(42, 8)),
	4203 => std_logic_vector(to_unsigned(42, 8)),
	4204 => std_logic_vector(to_unsigned(42, 8)),
	4205 => std_logic_vector(to_unsigned(41, 8)),
	4206 => std_logic_vector(to_unsigned(42, 8)),
	4207 => std_logic_vector(to_unsigned(41, 8)),
	4208 => std_logic_vector(to_unsigned(42, 8)),
	4209 => std_logic_vector(to_unsigned(42, 8)),
	4210 => std_logic_vector(to_unsigned(41, 8)),
	4211 => std_logic_vector(to_unsigned(41, 8)),
	4212 => std_logic_vector(to_unsigned(42, 8)),
	4213 => std_logic_vector(to_unsigned(42, 8)),
	4214 => std_logic_vector(to_unsigned(42, 8)),
	4215 => std_logic_vector(to_unsigned(42, 8)),
	4216 => std_logic_vector(to_unsigned(41, 8)),
	4217 => std_logic_vector(to_unsigned(41, 8)),
	4218 => std_logic_vector(to_unsigned(42, 8)),
	4219 => std_logic_vector(to_unsigned(42, 8)),
	4220 => std_logic_vector(to_unsigned(41, 8)),
	4221 => std_logic_vector(to_unsigned(42, 8)),
	4222 => std_logic_vector(to_unsigned(41, 8)),
	4223 => std_logic_vector(to_unsigned(42, 8)),
	4224 => std_logic_vector(to_unsigned(42, 8)),
	4225 => std_logic_vector(to_unsigned(41, 8)),
	4226 => std_logic_vector(to_unsigned(42, 8)),
	4227 => std_logic_vector(to_unsigned(41, 8)),
	4228 => std_logic_vector(to_unsigned(41, 8)),
	4229 => std_logic_vector(to_unsigned(41, 8)),
	4230 => std_logic_vector(to_unsigned(42, 8)),
	4231 => std_logic_vector(to_unsigned(41, 8)),
	4232 => std_logic_vector(to_unsigned(41, 8)),
	4233 => std_logic_vector(to_unsigned(41, 8)),
	4234 => std_logic_vector(to_unsigned(41, 8)),
	4235 => std_logic_vector(to_unsigned(41, 8)),
	4236 => std_logic_vector(to_unsigned(41, 8)),
	4237 => std_logic_vector(to_unsigned(41, 8)),
	4238 => std_logic_vector(to_unsigned(41, 8)),
	4239 => std_logic_vector(to_unsigned(42, 8)),
	4240 => std_logic_vector(to_unsigned(41, 8)),
	4241 => std_logic_vector(to_unsigned(42, 8)),
	4242 => std_logic_vector(to_unsigned(42, 8)),
	4243 => std_logic_vector(to_unsigned(42, 8)),
	4244 => std_logic_vector(to_unsigned(41, 8)),
	4245 => std_logic_vector(to_unsigned(41, 8)),
	4246 => std_logic_vector(to_unsigned(42, 8)),
	4247 => std_logic_vector(to_unsigned(41, 8)),
	4248 => std_logic_vector(to_unsigned(42, 8)),
	4249 => std_logic_vector(to_unsigned(41, 8)),
	4250 => std_logic_vector(to_unsigned(41, 8)),
	4251 => std_logic_vector(to_unsigned(41, 8)),
	4252 => std_logic_vector(to_unsigned(41, 8)),
	4253 => std_logic_vector(to_unsigned(41, 8)),
	4254 => std_logic_vector(to_unsigned(42, 8)),
	4255 => std_logic_vector(to_unsigned(42, 8)),
	4256 => std_logic_vector(to_unsigned(42, 8)),
	4257 => std_logic_vector(to_unsigned(41, 8)),
	4258 => std_logic_vector(to_unsigned(42, 8)),
	4259 => std_logic_vector(to_unsigned(42, 8)),
	4260 => std_logic_vector(to_unsigned(41, 8)),
	4261 => std_logic_vector(to_unsigned(41, 8)),
	4262 => std_logic_vector(to_unsigned(42, 8)),
	4263 => std_logic_vector(to_unsigned(42, 8)),
	4264 => std_logic_vector(to_unsigned(41, 8)),
	4265 => std_logic_vector(to_unsigned(41, 8)),
	4266 => std_logic_vector(to_unsigned(42, 8)),
	4267 => std_logic_vector(to_unsigned(41, 8)),
	4268 => std_logic_vector(to_unsigned(41, 8)),
	4269 => std_logic_vector(to_unsigned(41, 8)),
	4270 => std_logic_vector(to_unsigned(41, 8)),
	4271 => std_logic_vector(to_unsigned(41, 8)),
	4272 => std_logic_vector(to_unsigned(41, 8)),
	4273 => std_logic_vector(to_unsigned(41, 8)),
	4274 => std_logic_vector(to_unsigned(42, 8)),
	4275 => std_logic_vector(to_unsigned(42, 8)),
	4276 => std_logic_vector(to_unsigned(42, 8)),
	4277 => std_logic_vector(to_unsigned(41, 8)),
	4278 => std_logic_vector(to_unsigned(41, 8)),
	4279 => std_logic_vector(to_unsigned(42, 8)),
	4280 => std_logic_vector(to_unsigned(42, 8)),
	4281 => std_logic_vector(to_unsigned(41, 8)),
	4282 => std_logic_vector(to_unsigned(42, 8)),
	4283 => std_logic_vector(to_unsigned(42, 8)),
	4284 => std_logic_vector(to_unsigned(42, 8)),
	4285 => std_logic_vector(to_unsigned(42, 8)),
	4286 => std_logic_vector(to_unsigned(41, 8)),
	4287 => std_logic_vector(to_unsigned(42, 8)),
	4288 => std_logic_vector(to_unsigned(41, 8)),
	4289 => std_logic_vector(to_unsigned(41, 8)),
	4290 => std_logic_vector(to_unsigned(42, 8)),
	4291 => std_logic_vector(to_unsigned(42, 8)),
	4292 => std_logic_vector(to_unsigned(41, 8)),
	4293 => std_logic_vector(to_unsigned(41, 8)),
	4294 => std_logic_vector(to_unsigned(41, 8)),
	4295 => std_logic_vector(to_unsigned(41, 8)),
	4296 => std_logic_vector(to_unsigned(41, 8)),
	4297 => std_logic_vector(to_unsigned(42, 8)),
	4298 => std_logic_vector(to_unsigned(42, 8)),
	4299 => std_logic_vector(to_unsigned(41, 8)),
	4300 => std_logic_vector(to_unsigned(41, 8)),
	4301 => std_logic_vector(to_unsigned(42, 8)),
	4302 => std_logic_vector(to_unsigned(41, 8)),
	4303 => std_logic_vector(to_unsigned(41, 8)),
	4304 => std_logic_vector(to_unsigned(41, 8)),
	4305 => std_logic_vector(to_unsigned(41, 8)),
	4306 => std_logic_vector(to_unsigned(41, 8)),
	4307 => std_logic_vector(to_unsigned(42, 8)),
	4308 => std_logic_vector(to_unsigned(41, 8)),
	4309 => std_logic_vector(to_unsigned(41, 8)),
	4310 => std_logic_vector(to_unsigned(42, 8)),
	4311 => std_logic_vector(to_unsigned(41, 8)),
	4312 => std_logic_vector(to_unsigned(41, 8)),
	4313 => std_logic_vector(to_unsigned(42, 8)),
	4314 => std_logic_vector(to_unsigned(42, 8)),
	4315 => std_logic_vector(to_unsigned(42, 8)),
	4316 => std_logic_vector(to_unsigned(41, 8)),
	4317 => std_logic_vector(to_unsigned(41, 8)),
	4318 => std_logic_vector(to_unsigned(41, 8)),
	4319 => std_logic_vector(to_unsigned(41, 8)),
	4320 => std_logic_vector(to_unsigned(41, 8)),
	4321 => std_logic_vector(to_unsigned(41, 8)),
	4322 => std_logic_vector(to_unsigned(42, 8)),
	4323 => std_logic_vector(to_unsigned(42, 8)),
	4324 => std_logic_vector(to_unsigned(41, 8)),
	4325 => std_logic_vector(to_unsigned(42, 8)),
	4326 => std_logic_vector(to_unsigned(41, 8)),
	4327 => std_logic_vector(to_unsigned(42, 8)),
	4328 => std_logic_vector(to_unsigned(41, 8)),
	4329 => std_logic_vector(to_unsigned(42, 8)),
	4330 => std_logic_vector(to_unsigned(41, 8)),
	4331 => std_logic_vector(to_unsigned(41, 8)),
	4332 => std_logic_vector(to_unsigned(42, 8)),
	4333 => std_logic_vector(to_unsigned(41, 8)),
	4334 => std_logic_vector(to_unsigned(41, 8)),
	4335 => std_logic_vector(to_unsigned(42, 8)),
	4336 => std_logic_vector(to_unsigned(42, 8)),
	4337 => std_logic_vector(to_unsigned(42, 8)),
	4338 => std_logic_vector(to_unsigned(41, 8)),
	4339 => std_logic_vector(to_unsigned(42, 8)),
	4340 => std_logic_vector(to_unsigned(41, 8)),
	4341 => std_logic_vector(to_unsigned(42, 8)),
	4342 => std_logic_vector(to_unsigned(41, 8)),
	4343 => std_logic_vector(to_unsigned(42, 8)),
	4344 => std_logic_vector(to_unsigned(42, 8)),
	4345 => std_logic_vector(to_unsigned(42, 8)),
	4346 => std_logic_vector(to_unsigned(42, 8)),
	4347 => std_logic_vector(to_unsigned(41, 8)),
	4348 => std_logic_vector(to_unsigned(42, 8)),
	4349 => std_logic_vector(to_unsigned(41, 8)),
	4350 => std_logic_vector(to_unsigned(41, 8)),
	4351 => std_logic_vector(to_unsigned(41, 8)),
	4352 => std_logic_vector(to_unsigned(42, 8)),
	4353 => std_logic_vector(to_unsigned(42, 8)),
	4354 => std_logic_vector(to_unsigned(41, 8)),
	4355 => std_logic_vector(to_unsigned(41, 8)),
	4356 => std_logic_vector(to_unsigned(41, 8)),
	4357 => std_logic_vector(to_unsigned(42, 8)),
	4358 => std_logic_vector(to_unsigned(41, 8)),
	4359 => std_logic_vector(to_unsigned(41, 8)),
	4360 => std_logic_vector(to_unsigned(41, 8)),
	4361 => std_logic_vector(to_unsigned(42, 8)),
	4362 => std_logic_vector(to_unsigned(41, 8)),
	4363 => std_logic_vector(to_unsigned(42, 8)),
	4364 => std_logic_vector(to_unsigned(42, 8)),
	4365 => std_logic_vector(to_unsigned(42, 8)),
	4366 => std_logic_vector(to_unsigned(42, 8)),
	4367 => std_logic_vector(to_unsigned(42, 8)),
	4368 => std_logic_vector(to_unsigned(42, 8)),
	4369 => std_logic_vector(to_unsigned(41, 8)),
	4370 => std_logic_vector(to_unsigned(42, 8)),
	4371 => std_logic_vector(to_unsigned(41, 8)),
	4372 => std_logic_vector(to_unsigned(42, 8)),
	4373 => std_logic_vector(to_unsigned(41, 8)),
	4374 => std_logic_vector(to_unsigned(41, 8)),
	4375 => std_logic_vector(to_unsigned(41, 8)),
	4376 => std_logic_vector(to_unsigned(41, 8)),
	4377 => std_logic_vector(to_unsigned(42, 8)),
	4378 => std_logic_vector(to_unsigned(41, 8)),
	4379 => std_logic_vector(to_unsigned(41, 8)),
	4380 => std_logic_vector(to_unsigned(41, 8)),
	4381 => std_logic_vector(to_unsigned(41, 8)),
	4382 => std_logic_vector(to_unsigned(41, 8)),
	4383 => std_logic_vector(to_unsigned(41, 8)),
	4384 => std_logic_vector(to_unsigned(42, 8)),
	4385 => std_logic_vector(to_unsigned(41, 8)),
	4386 => std_logic_vector(to_unsigned(41, 8)),
	4387 => std_logic_vector(to_unsigned(42, 8)),
	4388 => std_logic_vector(to_unsigned(41, 8)),
	4389 => std_logic_vector(to_unsigned(42, 8)),
	4390 => std_logic_vector(to_unsigned(42, 8)),
	4391 => std_logic_vector(to_unsigned(42, 8)),
	4392 => std_logic_vector(to_unsigned(42, 8)),
	4393 => std_logic_vector(to_unsigned(41, 8)),
	4394 => std_logic_vector(to_unsigned(42, 8)),
	4395 => std_logic_vector(to_unsigned(41, 8)),
	4396 => std_logic_vector(to_unsigned(41, 8)),
	4397 => std_logic_vector(to_unsigned(41, 8)),
	4398 => std_logic_vector(to_unsigned(42, 8)),
	4399 => std_logic_vector(to_unsigned(42, 8)),
	4400 => std_logic_vector(to_unsigned(42, 8)),
	4401 => std_logic_vector(to_unsigned(41, 8)),
	4402 => std_logic_vector(to_unsigned(42, 8)),
	4403 => std_logic_vector(to_unsigned(42, 8)),
	4404 => std_logic_vector(to_unsigned(41, 8)),
	4405 => std_logic_vector(to_unsigned(42, 8)),
	4406 => std_logic_vector(to_unsigned(42, 8)),
	4407 => std_logic_vector(to_unsigned(42, 8)),
	4408 => std_logic_vector(to_unsigned(42, 8)),
	4409 => std_logic_vector(to_unsigned(41, 8)),
	4410 => std_logic_vector(to_unsigned(42, 8)),
	4411 => std_logic_vector(to_unsigned(42, 8)),
	4412 => std_logic_vector(to_unsigned(42, 8)),
	4413 => std_logic_vector(to_unsigned(42, 8)),
	4414 => std_logic_vector(to_unsigned(41, 8)),
	4415 => std_logic_vector(to_unsigned(42, 8)),
	4416 => std_logic_vector(to_unsigned(42, 8)),
	4417 => std_logic_vector(to_unsigned(41, 8)),
	4418 => std_logic_vector(to_unsigned(42, 8)),
	4419 => std_logic_vector(to_unsigned(41, 8)),
	4420 => std_logic_vector(to_unsigned(41, 8)),
	4421 => std_logic_vector(to_unsigned(42, 8)),
	4422 => std_logic_vector(to_unsigned(42, 8)),
	4423 => std_logic_vector(to_unsigned(41, 8)),
	4424 => std_logic_vector(to_unsigned(42, 8)),
	4425 => std_logic_vector(to_unsigned(41, 8)),
	4426 => std_logic_vector(to_unsigned(42, 8)),
	4427 => std_logic_vector(to_unsigned(41, 8)),
	4428 => std_logic_vector(to_unsigned(42, 8)),
	4429 => std_logic_vector(to_unsigned(42, 8)),
	4430 => std_logic_vector(to_unsigned(41, 8)),
	4431 => std_logic_vector(to_unsigned(41, 8)),
	4432 => std_logic_vector(to_unsigned(42, 8)),
	4433 => std_logic_vector(to_unsigned(41, 8)),
	4434 => std_logic_vector(to_unsigned(41, 8)),
	4435 => std_logic_vector(to_unsigned(41, 8)),
	4436 => std_logic_vector(to_unsigned(42, 8)),
	4437 => std_logic_vector(to_unsigned(42, 8)),
	4438 => std_logic_vector(to_unsigned(42, 8)),
	4439 => std_logic_vector(to_unsigned(41, 8)),
	4440 => std_logic_vector(to_unsigned(42, 8)),
	4441 => std_logic_vector(to_unsigned(41, 8)),
	4442 => std_logic_vector(to_unsigned(42, 8)),
	4443 => std_logic_vector(to_unsigned(42, 8)),
	4444 => std_logic_vector(to_unsigned(42, 8)),
	4445 => std_logic_vector(to_unsigned(41, 8)),
	4446 => std_logic_vector(to_unsigned(42, 8)),
	4447 => std_logic_vector(to_unsigned(41, 8)),
	4448 => std_logic_vector(to_unsigned(41, 8)),
	4449 => std_logic_vector(to_unsigned(41, 8)),
	4450 => std_logic_vector(to_unsigned(41, 8)),
	4451 => std_logic_vector(to_unsigned(42, 8)),
	4452 => std_logic_vector(to_unsigned(41, 8)),
	4453 => std_logic_vector(to_unsigned(42, 8)),
	4454 => std_logic_vector(to_unsigned(42, 8)),
	4455 => std_logic_vector(to_unsigned(42, 8)),
	4456 => std_logic_vector(to_unsigned(41, 8)),
	4457 => std_logic_vector(to_unsigned(42, 8)),
	4458 => std_logic_vector(to_unsigned(41, 8)),
	4459 => std_logic_vector(to_unsigned(41, 8)),
	4460 => std_logic_vector(to_unsigned(42, 8)),
	4461 => std_logic_vector(to_unsigned(41, 8)),
	4462 => std_logic_vector(to_unsigned(41, 8)),
	4463 => std_logic_vector(to_unsigned(41, 8)),
	4464 => std_logic_vector(to_unsigned(41, 8)),
	4465 => std_logic_vector(to_unsigned(41, 8)),
	4466 => std_logic_vector(to_unsigned(42, 8)),
	4467 => std_logic_vector(to_unsigned(42, 8)),
	4468 => std_logic_vector(to_unsigned(41, 8)),
	4469 => std_logic_vector(to_unsigned(42, 8)),
	4470 => std_logic_vector(to_unsigned(41, 8)),
	4471 => std_logic_vector(to_unsigned(42, 8)),
	4472 => std_logic_vector(to_unsigned(42, 8)),
	4473 => std_logic_vector(to_unsigned(41, 8)),
	4474 => std_logic_vector(to_unsigned(41, 8)),
	4475 => std_logic_vector(to_unsigned(42, 8)),
	4476 => std_logic_vector(to_unsigned(42, 8)),
	4477 => std_logic_vector(to_unsigned(42, 8)),
	4478 => std_logic_vector(to_unsigned(42, 8)),
	4479 => std_logic_vector(to_unsigned(42, 8)),
	4480 => std_logic_vector(to_unsigned(41, 8)),
	4481 => std_logic_vector(to_unsigned(41, 8)),
	4482 => std_logic_vector(to_unsigned(41, 8)),
	4483 => std_logic_vector(to_unsigned(42, 8)),
	4484 => std_logic_vector(to_unsigned(41, 8)),
	4485 => std_logic_vector(to_unsigned(41, 8)),
	4486 => std_logic_vector(to_unsigned(42, 8)),
	4487 => std_logic_vector(to_unsigned(42, 8)),
	4488 => std_logic_vector(to_unsigned(42, 8)),
	4489 => std_logic_vector(to_unsigned(41, 8)),
	4490 => std_logic_vector(to_unsigned(41, 8)),
	4491 => std_logic_vector(to_unsigned(41, 8)),
	4492 => std_logic_vector(to_unsigned(42, 8)),
	4493 => std_logic_vector(to_unsigned(41, 8)),
	4494 => std_logic_vector(to_unsigned(41, 8)),
	4495 => std_logic_vector(to_unsigned(42, 8)),
	4496 => std_logic_vector(to_unsigned(41, 8)),
	4497 => std_logic_vector(to_unsigned(42, 8)),
	4498 => std_logic_vector(to_unsigned(41, 8)),
	4499 => std_logic_vector(to_unsigned(42, 8)),
	4500 => std_logic_vector(to_unsigned(42, 8)),
	4501 => std_logic_vector(to_unsigned(41, 8)),
	4502 => std_logic_vector(to_unsigned(42, 8)),
	4503 => std_logic_vector(to_unsigned(42, 8)),
	4504 => std_logic_vector(to_unsigned(41, 8)),
	4505 => std_logic_vector(to_unsigned(41, 8)),
	4506 => std_logic_vector(to_unsigned(41, 8)),
	4507 => std_logic_vector(to_unsigned(42, 8)),
	4508 => std_logic_vector(to_unsigned(41, 8)),
	4509 => std_logic_vector(to_unsigned(42, 8)),
	4510 => std_logic_vector(to_unsigned(42, 8)),
	4511 => std_logic_vector(to_unsigned(41, 8)),
	4512 => std_logic_vector(to_unsigned(41, 8)),
	4513 => std_logic_vector(to_unsigned(41, 8)),
	4514 => std_logic_vector(to_unsigned(41, 8)),
	4515 => std_logic_vector(to_unsigned(42, 8)),
	4516 => std_logic_vector(to_unsigned(42, 8)),
	4517 => std_logic_vector(to_unsigned(42, 8)),
	4518 => std_logic_vector(to_unsigned(41, 8)),
	4519 => std_logic_vector(to_unsigned(41, 8)),
	4520 => std_logic_vector(to_unsigned(42, 8)),
	4521 => std_logic_vector(to_unsigned(42, 8)),
	4522 => std_logic_vector(to_unsigned(41, 8)),
	4523 => std_logic_vector(to_unsigned(41, 8)),
	4524 => std_logic_vector(to_unsigned(41, 8)),
	4525 => std_logic_vector(to_unsigned(41, 8)),
	4526 => std_logic_vector(to_unsigned(41, 8)),
	4527 => std_logic_vector(to_unsigned(41, 8)),
	4528 => std_logic_vector(to_unsigned(41, 8)),
	4529 => std_logic_vector(to_unsigned(41, 8)),
	4530 => std_logic_vector(to_unsigned(42, 8)),
	4531 => std_logic_vector(to_unsigned(41, 8)),
	4532 => std_logic_vector(to_unsigned(41, 8)),
	4533 => std_logic_vector(to_unsigned(41, 8)),
	4534 => std_logic_vector(to_unsigned(41, 8)),
	4535 => std_logic_vector(to_unsigned(42, 8)),
	4536 => std_logic_vector(to_unsigned(42, 8)),
	4537 => std_logic_vector(to_unsigned(42, 8)),
	4538 => std_logic_vector(to_unsigned(41, 8)),
	4539 => std_logic_vector(to_unsigned(41, 8)),
	4540 => std_logic_vector(to_unsigned(42, 8)),
	4541 => std_logic_vector(to_unsigned(42, 8)),
	4542 => std_logic_vector(to_unsigned(42, 8)),
	4543 => std_logic_vector(to_unsigned(41, 8)),
	4544 => std_logic_vector(to_unsigned(41, 8)),
	4545 => std_logic_vector(to_unsigned(41, 8)),
	4546 => std_logic_vector(to_unsigned(42, 8)),
	4547 => std_logic_vector(to_unsigned(42, 8)),
	4548 => std_logic_vector(to_unsigned(42, 8)),
	4549 => std_logic_vector(to_unsigned(41, 8)),
	4550 => std_logic_vector(to_unsigned(41, 8)),
	4551 => std_logic_vector(to_unsigned(41, 8)),
	4552 => std_logic_vector(to_unsigned(41, 8)),
	4553 => std_logic_vector(to_unsigned(41, 8)),
	4554 => std_logic_vector(to_unsigned(41, 8)),
	4555 => std_logic_vector(to_unsigned(41, 8)),
	4556 => std_logic_vector(to_unsigned(42, 8)),
	4557 => std_logic_vector(to_unsigned(41, 8)),
	4558 => std_logic_vector(to_unsigned(41, 8)),
	4559 => std_logic_vector(to_unsigned(42, 8)),
	4560 => std_logic_vector(to_unsigned(41, 8)),
	4561 => std_logic_vector(to_unsigned(41, 8)),
	4562 => std_logic_vector(to_unsigned(41, 8)),
	4563 => std_logic_vector(to_unsigned(41, 8)),
	4564 => std_logic_vector(to_unsigned(41, 8)),
	4565 => std_logic_vector(to_unsigned(42, 8)),
	4566 => std_logic_vector(to_unsigned(41, 8)),
	4567 => std_logic_vector(to_unsigned(41, 8)),
	4568 => std_logic_vector(to_unsigned(42, 8)),
	4569 => std_logic_vector(to_unsigned(41, 8)),
	4570 => std_logic_vector(to_unsigned(42, 8)),
	4571 => std_logic_vector(to_unsigned(41, 8)),
	4572 => std_logic_vector(to_unsigned(41, 8)),
	4573 => std_logic_vector(to_unsigned(41, 8)),
	4574 => std_logic_vector(to_unsigned(41, 8)),
	4575 => std_logic_vector(to_unsigned(42, 8)),
	4576 => std_logic_vector(to_unsigned(41, 8)),
	4577 => std_logic_vector(to_unsigned(42, 8)),
	4578 => std_logic_vector(to_unsigned(41, 8)),
	4579 => std_logic_vector(to_unsigned(41, 8)),
	4580 => std_logic_vector(to_unsigned(41, 8)),
	4581 => std_logic_vector(to_unsigned(42, 8)),
	4582 => std_logic_vector(to_unsigned(42, 8)),
	4583 => std_logic_vector(to_unsigned(42, 8)),
	4584 => std_logic_vector(to_unsigned(41, 8)),
	4585 => std_logic_vector(to_unsigned(42, 8)),
	4586 => std_logic_vector(to_unsigned(41, 8)),
	4587 => std_logic_vector(to_unsigned(42, 8)),
	4588 => std_logic_vector(to_unsigned(41, 8)),
	4589 => std_logic_vector(to_unsigned(41, 8)),
	4590 => std_logic_vector(to_unsigned(42, 8)),
	4591 => std_logic_vector(to_unsigned(42, 8)),
	4592 => std_logic_vector(to_unsigned(42, 8)),
	4593 => std_logic_vector(to_unsigned(42, 8)),
	4594 => std_logic_vector(to_unsigned(41, 8)),
	4595 => std_logic_vector(to_unsigned(42, 8)),
	4596 => std_logic_vector(to_unsigned(41, 8)),
	4597 => std_logic_vector(to_unsigned(41, 8)),
	4598 => std_logic_vector(to_unsigned(42, 8)),
	4599 => std_logic_vector(to_unsigned(42, 8)),
	4600 => std_logic_vector(to_unsigned(42, 8)),
	4601 => std_logic_vector(to_unsigned(42, 8)),
	4602 => std_logic_vector(to_unsigned(42, 8)),
	4603 => std_logic_vector(to_unsigned(42, 8)),
	4604 => std_logic_vector(to_unsigned(42, 8)),
	4605 => std_logic_vector(to_unsigned(42, 8)),
	4606 => std_logic_vector(to_unsigned(41, 8)),
	4607 => std_logic_vector(to_unsigned(41, 8)),
	4608 => std_logic_vector(to_unsigned(41, 8)),
	4609 => std_logic_vector(to_unsigned(41, 8)),
	4610 => std_logic_vector(to_unsigned(42, 8)),
	4611 => std_logic_vector(to_unsigned(42, 8)),
	4612 => std_logic_vector(to_unsigned(42, 8)),
	4613 => std_logic_vector(to_unsigned(42, 8)),
	4614 => std_logic_vector(to_unsigned(42, 8)),
	4615 => std_logic_vector(to_unsigned(41, 8)),
	4616 => std_logic_vector(to_unsigned(41, 8)),
	4617 => std_logic_vector(to_unsigned(41, 8)),
	4618 => std_logic_vector(to_unsigned(41, 8)),
	4619 => std_logic_vector(to_unsigned(42, 8)),
	4620 => std_logic_vector(to_unsigned(42, 8)),
	4621 => std_logic_vector(to_unsigned(41, 8)),
	4622 => std_logic_vector(to_unsigned(42, 8)),
	4623 => std_logic_vector(to_unsigned(41, 8)),
	4624 => std_logic_vector(to_unsigned(41, 8)),
	4625 => std_logic_vector(to_unsigned(42, 8)),
	4626 => std_logic_vector(to_unsigned(41, 8)),
	4627 => std_logic_vector(to_unsigned(42, 8)),
	4628 => std_logic_vector(to_unsigned(42, 8)),
	4629 => std_logic_vector(to_unsigned(42, 8)),
	4630 => std_logic_vector(to_unsigned(42, 8)),
	4631 => std_logic_vector(to_unsigned(41, 8)),
	4632 => std_logic_vector(to_unsigned(41, 8)),
	4633 => std_logic_vector(to_unsigned(42, 8)),
	4634 => std_logic_vector(to_unsigned(42, 8)),
	4635 => std_logic_vector(to_unsigned(42, 8)),
	4636 => std_logic_vector(to_unsigned(42, 8)),
	4637 => std_logic_vector(to_unsigned(42, 8)),
	4638 => std_logic_vector(to_unsigned(41, 8)),
	4639 => std_logic_vector(to_unsigned(41, 8)),
	4640 => std_logic_vector(to_unsigned(41, 8)),
	4641 => std_logic_vector(to_unsigned(42, 8)),
	4642 => std_logic_vector(to_unsigned(42, 8)),
	4643 => std_logic_vector(to_unsigned(42, 8)),
	4644 => std_logic_vector(to_unsigned(41, 8)),
	4645 => std_logic_vector(to_unsigned(42, 8)),
	4646 => std_logic_vector(to_unsigned(42, 8)),
	4647 => std_logic_vector(to_unsigned(42, 8)),
	4648 => std_logic_vector(to_unsigned(41, 8)),
	4649 => std_logic_vector(to_unsigned(42, 8)),
	4650 => std_logic_vector(to_unsigned(42, 8)),
	4651 => std_logic_vector(to_unsigned(42, 8)),
	4652 => std_logic_vector(to_unsigned(41, 8)),
	4653 => std_logic_vector(to_unsigned(41, 8)),
	4654 => std_logic_vector(to_unsigned(42, 8)),
	4655 => std_logic_vector(to_unsigned(41, 8)),
	4656 => std_logic_vector(to_unsigned(41, 8)),
	4657 => std_logic_vector(to_unsigned(42, 8)),
	4658 => std_logic_vector(to_unsigned(42, 8)),
	4659 => std_logic_vector(to_unsigned(41, 8)),
	4660 => std_logic_vector(to_unsigned(41, 8)),
	4661 => std_logic_vector(to_unsigned(41, 8)),
	4662 => std_logic_vector(to_unsigned(42, 8)),
	4663 => std_logic_vector(to_unsigned(41, 8)),
	4664 => std_logic_vector(to_unsigned(41, 8)),
	4665 => std_logic_vector(to_unsigned(42, 8)),
	4666 => std_logic_vector(to_unsigned(41, 8)),
	4667 => std_logic_vector(to_unsigned(42, 8)),
	4668 => std_logic_vector(to_unsigned(42, 8)),
	4669 => std_logic_vector(to_unsigned(42, 8)),
	4670 => std_logic_vector(to_unsigned(42, 8)),
	4671 => std_logic_vector(to_unsigned(41, 8)),
	4672 => std_logic_vector(to_unsigned(42, 8)),
	4673 => std_logic_vector(to_unsigned(42, 8)),
	4674 => std_logic_vector(to_unsigned(42, 8)),
	4675 => std_logic_vector(to_unsigned(41, 8)),
	4676 => std_logic_vector(to_unsigned(42, 8)),
	4677 => std_logic_vector(to_unsigned(42, 8)),
	4678 => std_logic_vector(to_unsigned(42, 8)),
	4679 => std_logic_vector(to_unsigned(41, 8)),
	4680 => std_logic_vector(to_unsigned(42, 8)),
	4681 => std_logic_vector(to_unsigned(42, 8)),
	4682 => std_logic_vector(to_unsigned(42, 8)),
	4683 => std_logic_vector(to_unsigned(41, 8)),
	4684 => std_logic_vector(to_unsigned(42, 8)),
	4685 => std_logic_vector(to_unsigned(41, 8)),
	4686 => std_logic_vector(to_unsigned(42, 8)),
	4687 => std_logic_vector(to_unsigned(41, 8)),
	4688 => std_logic_vector(to_unsigned(42, 8)),
	4689 => std_logic_vector(to_unsigned(42, 8)),
	4690 => std_logic_vector(to_unsigned(42, 8)),
	4691 => std_logic_vector(to_unsigned(41, 8)),
	4692 => std_logic_vector(to_unsigned(42, 8)),
	4693 => std_logic_vector(to_unsigned(41, 8)),
	4694 => std_logic_vector(to_unsigned(42, 8)),
	4695 => std_logic_vector(to_unsigned(42, 8)),
	4696 => std_logic_vector(to_unsigned(42, 8)),
	4697 => std_logic_vector(to_unsigned(42, 8)),
	4698 => std_logic_vector(to_unsigned(42, 8)),
	4699 => std_logic_vector(to_unsigned(42, 8)),
	4700 => std_logic_vector(to_unsigned(42, 8)),
	4701 => std_logic_vector(to_unsigned(42, 8)),
	4702 => std_logic_vector(to_unsigned(42, 8)),
	4703 => std_logic_vector(to_unsigned(42, 8)),
	4704 => std_logic_vector(to_unsigned(41, 8)),
	4705 => std_logic_vector(to_unsigned(41, 8)),
	4706 => std_logic_vector(to_unsigned(42, 8)),
	4707 => std_logic_vector(to_unsigned(41, 8)),
	4708 => std_logic_vector(to_unsigned(41, 8)),
	4709 => std_logic_vector(to_unsigned(41, 8)),
	4710 => std_logic_vector(to_unsigned(41, 8)),
	4711 => std_logic_vector(to_unsigned(41, 8)),
	4712 => std_logic_vector(to_unsigned(41, 8)),
	4713 => std_logic_vector(to_unsigned(42, 8)),
	4714 => std_logic_vector(to_unsigned(42, 8)),
	4715 => std_logic_vector(to_unsigned(41, 8)),
	4716 => std_logic_vector(to_unsigned(42, 8)),
	4717 => std_logic_vector(to_unsigned(41, 8)),
	4718 => std_logic_vector(to_unsigned(42, 8)),
	4719 => std_logic_vector(to_unsigned(42, 8)),
	4720 => std_logic_vector(to_unsigned(42, 8)),
	4721 => std_logic_vector(to_unsigned(41, 8)),
	4722 => std_logic_vector(to_unsigned(41, 8)),
	4723 => std_logic_vector(to_unsigned(42, 8)),
	4724 => std_logic_vector(to_unsigned(42, 8)),
	4725 => std_logic_vector(to_unsigned(41, 8)),
	4726 => std_logic_vector(to_unsigned(42, 8)),
	4727 => std_logic_vector(to_unsigned(41, 8)),
	4728 => std_logic_vector(to_unsigned(41, 8)),
	4729 => std_logic_vector(to_unsigned(42, 8)),
	4730 => std_logic_vector(to_unsigned(42, 8)),
	4731 => std_logic_vector(to_unsigned(41, 8)),
	4732 => std_logic_vector(to_unsigned(41, 8)),
	4733 => std_logic_vector(to_unsigned(41, 8)),
	4734 => std_logic_vector(to_unsigned(41, 8)),
	4735 => std_logic_vector(to_unsigned(42, 8)),
	4736 => std_logic_vector(to_unsigned(41, 8)),
	4737 => std_logic_vector(to_unsigned(42, 8)),
	4738 => std_logic_vector(to_unsigned(42, 8)),
	4739 => std_logic_vector(to_unsigned(41, 8)),
	4740 => std_logic_vector(to_unsigned(41, 8)),
	4741 => std_logic_vector(to_unsigned(42, 8)),
	4742 => std_logic_vector(to_unsigned(41, 8)),
	4743 => std_logic_vector(to_unsigned(42, 8)),
	4744 => std_logic_vector(to_unsigned(41, 8)),
	4745 => std_logic_vector(to_unsigned(42, 8)),
	4746 => std_logic_vector(to_unsigned(41, 8)),
	4747 => std_logic_vector(to_unsigned(41, 8)),
	4748 => std_logic_vector(to_unsigned(41, 8)),
	4749 => std_logic_vector(to_unsigned(41, 8)),
	4750 => std_logic_vector(to_unsigned(41, 8)),
	4751 => std_logic_vector(to_unsigned(42, 8)),
	4752 => std_logic_vector(to_unsigned(41, 8)),
	4753 => std_logic_vector(to_unsigned(42, 8)),
	4754 => std_logic_vector(to_unsigned(42, 8)),
	4755 => std_logic_vector(to_unsigned(42, 8)),
	4756 => std_logic_vector(to_unsigned(42, 8)),
	4757 => std_logic_vector(to_unsigned(42, 8)),
	4758 => std_logic_vector(to_unsigned(42, 8)),
	4759 => std_logic_vector(to_unsigned(42, 8)),
	4760 => std_logic_vector(to_unsigned(42, 8)),
	4761 => std_logic_vector(to_unsigned(42, 8)),
	4762 => std_logic_vector(to_unsigned(41, 8)),
	4763 => std_logic_vector(to_unsigned(42, 8)),
	4764 => std_logic_vector(to_unsigned(41, 8)),
	4765 => std_logic_vector(to_unsigned(42, 8)),
	4766 => std_logic_vector(to_unsigned(41, 8)),
	4767 => std_logic_vector(to_unsigned(42, 8)),
	4768 => std_logic_vector(to_unsigned(42, 8)),
	4769 => std_logic_vector(to_unsigned(42, 8)),
	4770 => std_logic_vector(to_unsigned(42, 8)),
	4771 => std_logic_vector(to_unsigned(42, 8)),
	4772 => std_logic_vector(to_unsigned(42, 8)),
	4773 => std_logic_vector(to_unsigned(41, 8)),
	4774 => std_logic_vector(to_unsigned(42, 8)),
	4775 => std_logic_vector(to_unsigned(42, 8)),
	4776 => std_logic_vector(to_unsigned(42, 8)),
	4777 => std_logic_vector(to_unsigned(41, 8)),
	4778 => std_logic_vector(to_unsigned(42, 8)),
	4779 => std_logic_vector(to_unsigned(41, 8)),
	4780 => std_logic_vector(to_unsigned(42, 8)),
	4781 => std_logic_vector(to_unsigned(42, 8)),
	4782 => std_logic_vector(to_unsigned(41, 8)),
	4783 => std_logic_vector(to_unsigned(41, 8)),
	4784 => std_logic_vector(to_unsigned(42, 8)),
	4785 => std_logic_vector(to_unsigned(41, 8)),
	4786 => std_logic_vector(to_unsigned(41, 8)),
	4787 => std_logic_vector(to_unsigned(42, 8)),
	4788 => std_logic_vector(to_unsigned(42, 8)),
	4789 => std_logic_vector(to_unsigned(42, 8)),
	4790 => std_logic_vector(to_unsigned(42, 8)),
	4791 => std_logic_vector(to_unsigned(41, 8)),
	4792 => std_logic_vector(to_unsigned(42, 8)),
	4793 => std_logic_vector(to_unsigned(42, 8)),
	4794 => std_logic_vector(to_unsigned(41, 8)),
	4795 => std_logic_vector(to_unsigned(41, 8)),
	4796 => std_logic_vector(to_unsigned(41, 8)),
	4797 => std_logic_vector(to_unsigned(41, 8)),
	4798 => std_logic_vector(to_unsigned(41, 8)),
	4799 => std_logic_vector(to_unsigned(41, 8)),
	4800 => std_logic_vector(to_unsigned(41, 8)),
	4801 => std_logic_vector(to_unsigned(42, 8)),
	4802 => std_logic_vector(to_unsigned(42, 8)),
	4803 => std_logic_vector(to_unsigned(42, 8)),
	4804 => std_logic_vector(to_unsigned(41, 8)),
	4805 => std_logic_vector(to_unsigned(41, 8)),
	4806 => std_logic_vector(to_unsigned(42, 8)),
	4807 => std_logic_vector(to_unsigned(42, 8)),
	4808 => std_logic_vector(to_unsigned(41, 8)),
	4809 => std_logic_vector(to_unsigned(41, 8)),
	4810 => std_logic_vector(to_unsigned(42, 8)),
	4811 => std_logic_vector(to_unsigned(41, 8)),
	4812 => std_logic_vector(to_unsigned(41, 8)),
	4813 => std_logic_vector(to_unsigned(42, 8)),
	4814 => std_logic_vector(to_unsigned(42, 8)),
	4815 => std_logic_vector(to_unsigned(42, 8)),
	4816 => std_logic_vector(to_unsigned(42, 8)),
	4817 => std_logic_vector(to_unsigned(42, 8)),
	4818 => std_logic_vector(to_unsigned(41, 8)),
	4819 => std_logic_vector(to_unsigned(41, 8)),
	4820 => std_logic_vector(to_unsigned(41, 8)),
	4821 => std_logic_vector(to_unsigned(42, 8)),
	4822 => std_logic_vector(to_unsigned(42, 8)),
	4823 => std_logic_vector(to_unsigned(42, 8)),
	4824 => std_logic_vector(to_unsigned(42, 8)),
	4825 => std_logic_vector(to_unsigned(42, 8)),
	4826 => std_logic_vector(to_unsigned(41, 8)),
	4827 => std_logic_vector(to_unsigned(42, 8)),
	4828 => std_logic_vector(to_unsigned(41, 8)),
	4829 => std_logic_vector(to_unsigned(42, 8)),
	4830 => std_logic_vector(to_unsigned(41, 8)),
	4831 => std_logic_vector(to_unsigned(41, 8)),
	4832 => std_logic_vector(to_unsigned(42, 8)),
	4833 => std_logic_vector(to_unsigned(42, 8)),
	4834 => std_logic_vector(to_unsigned(41, 8)),
	4835 => std_logic_vector(to_unsigned(42, 8)),
	4836 => std_logic_vector(to_unsigned(42, 8)),
	4837 => std_logic_vector(to_unsigned(41, 8)),
	4838 => std_logic_vector(to_unsigned(41, 8)),
	4839 => std_logic_vector(to_unsigned(42, 8)),
	4840 => std_logic_vector(to_unsigned(42, 8)),
	4841 => std_logic_vector(to_unsigned(41, 8)),
	4842 => std_logic_vector(to_unsigned(41, 8)),
	4843 => std_logic_vector(to_unsigned(41, 8)),
	4844 => std_logic_vector(to_unsigned(41, 8)),
	4845 => std_logic_vector(to_unsigned(41, 8)),
	4846 => std_logic_vector(to_unsigned(41, 8)),
	4847 => std_logic_vector(to_unsigned(41, 8)),
	4848 => std_logic_vector(to_unsigned(42, 8)),
	4849 => std_logic_vector(to_unsigned(41, 8)),
	4850 => std_logic_vector(to_unsigned(41, 8)),
	4851 => std_logic_vector(to_unsigned(42, 8)),
	4852 => std_logic_vector(to_unsigned(41, 8)),
	4853 => std_logic_vector(to_unsigned(42, 8)),
	4854 => std_logic_vector(to_unsigned(42, 8)),
	4855 => std_logic_vector(to_unsigned(41, 8)),
	4856 => std_logic_vector(to_unsigned(42, 8)),
	4857 => std_logic_vector(to_unsigned(41, 8)),
	4858 => std_logic_vector(to_unsigned(41, 8)),
	4859 => std_logic_vector(to_unsigned(41, 8)),
	4860 => std_logic_vector(to_unsigned(42, 8)),
	4861 => std_logic_vector(to_unsigned(42, 8)),
	4862 => std_logic_vector(to_unsigned(41, 8)),
	4863 => std_logic_vector(to_unsigned(42, 8)),
	4864 => std_logic_vector(to_unsigned(42, 8)),
	4865 => std_logic_vector(to_unsigned(41, 8)),
	4866 => std_logic_vector(to_unsigned(41, 8)),
	4867 => std_logic_vector(to_unsigned(42, 8)),
	4868 => std_logic_vector(to_unsigned(42, 8)),
	4869 => std_logic_vector(to_unsigned(42, 8)),
	4870 => std_logic_vector(to_unsigned(42, 8)),
	4871 => std_logic_vector(to_unsigned(41, 8)),
	4872 => std_logic_vector(to_unsigned(42, 8)),
	4873 => std_logic_vector(to_unsigned(41, 8)),
	4874 => std_logic_vector(to_unsigned(41, 8)),
	4875 => std_logic_vector(to_unsigned(42, 8)),
	4876 => std_logic_vector(to_unsigned(42, 8)),
	4877 => std_logic_vector(to_unsigned(41, 8)),
	4878 => std_logic_vector(to_unsigned(42, 8)),
	4879 => std_logic_vector(to_unsigned(42, 8)),
	4880 => std_logic_vector(to_unsigned(42, 8)),
	4881 => std_logic_vector(to_unsigned(42, 8)),
	4882 => std_logic_vector(to_unsigned(42, 8)),
	4883 => std_logic_vector(to_unsigned(41, 8)),
	4884 => std_logic_vector(to_unsigned(42, 8)),
	4885 => std_logic_vector(to_unsigned(41, 8)),
	4886 => std_logic_vector(to_unsigned(42, 8)),
	4887 => std_logic_vector(to_unsigned(41, 8)),
	4888 => std_logic_vector(to_unsigned(41, 8)),
	4889 => std_logic_vector(to_unsigned(41, 8)),
	4890 => std_logic_vector(to_unsigned(41, 8)),
	4891 => std_logic_vector(to_unsigned(42, 8)),
	4892 => std_logic_vector(to_unsigned(41, 8)),
	4893 => std_logic_vector(to_unsigned(41, 8)),
	4894 => std_logic_vector(to_unsigned(41, 8)),
	4895 => std_logic_vector(to_unsigned(42, 8)),
	4896 => std_logic_vector(to_unsigned(42, 8)),
	4897 => std_logic_vector(to_unsigned(41, 8)),
	4898 => std_logic_vector(to_unsigned(42, 8)),
	4899 => std_logic_vector(to_unsigned(41, 8)),
	4900 => std_logic_vector(to_unsigned(42, 8)),
	4901 => std_logic_vector(to_unsigned(42, 8)),
	4902 => std_logic_vector(to_unsigned(42, 8)),
	4903 => std_logic_vector(to_unsigned(42, 8)),
	4904 => std_logic_vector(to_unsigned(41, 8)),
	4905 => std_logic_vector(to_unsigned(41, 8)),
	4906 => std_logic_vector(to_unsigned(42, 8)),
	4907 => std_logic_vector(to_unsigned(42, 8)),
	4908 => std_logic_vector(to_unsigned(42, 8)),
	4909 => std_logic_vector(to_unsigned(42, 8)),
	4910 => std_logic_vector(to_unsigned(42, 8)),
	4911 => std_logic_vector(to_unsigned(41, 8)),
	4912 => std_logic_vector(to_unsigned(41, 8)),
	4913 => std_logic_vector(to_unsigned(42, 8)),
	4914 => std_logic_vector(to_unsigned(42, 8)),
	4915 => std_logic_vector(to_unsigned(41, 8)),
	4916 => std_logic_vector(to_unsigned(41, 8)),
	4917 => std_logic_vector(to_unsigned(42, 8)),
	4918 => std_logic_vector(to_unsigned(42, 8)),
	4919 => std_logic_vector(to_unsigned(41, 8)),
	4920 => std_logic_vector(to_unsigned(41, 8)),
	4921 => std_logic_vector(to_unsigned(42, 8)),
	4922 => std_logic_vector(to_unsigned(41, 8)),
	4923 => std_logic_vector(to_unsigned(41, 8)),
	4924 => std_logic_vector(to_unsigned(42, 8)),
	4925 => std_logic_vector(to_unsigned(42, 8)),
	4926 => std_logic_vector(to_unsigned(41, 8)),
	4927 => std_logic_vector(to_unsigned(41, 8)),
	4928 => std_logic_vector(to_unsigned(41, 8)),
	4929 => std_logic_vector(to_unsigned(42, 8)),
	4930 => std_logic_vector(to_unsigned(42, 8)),
	4931 => std_logic_vector(to_unsigned(41, 8)),
	4932 => std_logic_vector(to_unsigned(42, 8)),
	4933 => std_logic_vector(to_unsigned(41, 8)),
	4934 => std_logic_vector(to_unsigned(41, 8)),
	4935 => std_logic_vector(to_unsigned(41, 8)),
	4936 => std_logic_vector(to_unsigned(42, 8)),
	4937 => std_logic_vector(to_unsigned(41, 8)),
	4938 => std_logic_vector(to_unsigned(42, 8)),
	4939 => std_logic_vector(to_unsigned(41, 8)),
	4940 => std_logic_vector(to_unsigned(42, 8)),
	4941 => std_logic_vector(to_unsigned(42, 8)),
	4942 => std_logic_vector(to_unsigned(42, 8)),
	4943 => std_logic_vector(to_unsigned(42, 8)),
	4944 => std_logic_vector(to_unsigned(41, 8)),
	4945 => std_logic_vector(to_unsigned(42, 8)),
	4946 => std_logic_vector(to_unsigned(41, 8)),
	4947 => std_logic_vector(to_unsigned(42, 8)),
	4948 => std_logic_vector(to_unsigned(41, 8)),
	4949 => std_logic_vector(to_unsigned(41, 8)),
	4950 => std_logic_vector(to_unsigned(41, 8)),
	4951 => std_logic_vector(to_unsigned(42, 8)),
	4952 => std_logic_vector(to_unsigned(41, 8)),
	4953 => std_logic_vector(to_unsigned(41, 8)),
	4954 => std_logic_vector(to_unsigned(42, 8)),
	4955 => std_logic_vector(to_unsigned(42, 8)),
	4956 => std_logic_vector(to_unsigned(41, 8)),
	4957 => std_logic_vector(to_unsigned(41, 8)),
	4958 => std_logic_vector(to_unsigned(41, 8)),
	4959 => std_logic_vector(to_unsigned(42, 8)),
	4960 => std_logic_vector(to_unsigned(41, 8)),
	4961 => std_logic_vector(to_unsigned(42, 8)),
	4962 => std_logic_vector(to_unsigned(41, 8)),
	4963 => std_logic_vector(to_unsigned(41, 8)),
	4964 => std_logic_vector(to_unsigned(41, 8)),
	4965 => std_logic_vector(to_unsigned(41, 8)),
	4966 => std_logic_vector(to_unsigned(42, 8)),
	4967 => std_logic_vector(to_unsigned(41, 8)),
	4968 => std_logic_vector(to_unsigned(41, 8)),
	4969 => std_logic_vector(to_unsigned(42, 8)),
	4970 => std_logic_vector(to_unsigned(42, 8)),
	4971 => std_logic_vector(to_unsigned(42, 8)),
	4972 => std_logic_vector(to_unsigned(41, 8)),
	4973 => std_logic_vector(to_unsigned(42, 8)),
	4974 => std_logic_vector(to_unsigned(41, 8)),
	4975 => std_logic_vector(to_unsigned(42, 8)),
	4976 => std_logic_vector(to_unsigned(41, 8)),
	4977 => std_logic_vector(to_unsigned(41, 8)),
	4978 => std_logic_vector(to_unsigned(42, 8)),
	4979 => std_logic_vector(to_unsigned(42, 8)),
	4980 => std_logic_vector(to_unsigned(41, 8)),
	4981 => std_logic_vector(to_unsigned(41, 8)),
	4982 => std_logic_vector(to_unsigned(41, 8)),
	4983 => std_logic_vector(to_unsigned(42, 8)),
	4984 => std_logic_vector(to_unsigned(42, 8)),
	4985 => std_logic_vector(to_unsigned(42, 8)),
	4986 => std_logic_vector(to_unsigned(42, 8)),
	4987 => std_logic_vector(to_unsigned(42, 8)),
	4988 => std_logic_vector(to_unsigned(42, 8)),
	4989 => std_logic_vector(to_unsigned(41, 8)),
	4990 => std_logic_vector(to_unsigned(42, 8)),
	4991 => std_logic_vector(to_unsigned(41, 8)),
	4992 => std_logic_vector(to_unsigned(41, 8)),
	4993 => std_logic_vector(to_unsigned(42, 8)),
	4994 => std_logic_vector(to_unsigned(41, 8)),
	4995 => std_logic_vector(to_unsigned(41, 8)),
	4996 => std_logic_vector(to_unsigned(42, 8)),
	4997 => std_logic_vector(to_unsigned(42, 8)),
	4998 => std_logic_vector(to_unsigned(42, 8)),
	4999 => std_logic_vector(to_unsigned(42, 8)),
	5000 => std_logic_vector(to_unsigned(41, 8)),
	5001 => std_logic_vector(to_unsigned(42, 8)),
	5002 => std_logic_vector(to_unsigned(42, 8)),
	5003 => std_logic_vector(to_unsigned(41, 8)),
	5004 => std_logic_vector(to_unsigned(42, 8)),
	5005 => std_logic_vector(to_unsigned(41, 8)),
	5006 => std_logic_vector(to_unsigned(42, 8)),
	5007 => std_logic_vector(to_unsigned(41, 8)),
	5008 => std_logic_vector(to_unsigned(42, 8)),
	5009 => std_logic_vector(to_unsigned(41, 8)),
	5010 => std_logic_vector(to_unsigned(42, 8)),
	5011 => std_logic_vector(to_unsigned(42, 8)),
	5012 => std_logic_vector(to_unsigned(42, 8)),
	5013 => std_logic_vector(to_unsigned(41, 8)),
	5014 => std_logic_vector(to_unsigned(42, 8)),
	5015 => std_logic_vector(to_unsigned(41, 8)),
	5016 => std_logic_vector(to_unsigned(42, 8)),
	5017 => std_logic_vector(to_unsigned(41, 8)),
	5018 => std_logic_vector(to_unsigned(41, 8)),
	5019 => std_logic_vector(to_unsigned(42, 8)),
	5020 => std_logic_vector(to_unsigned(42, 8)),
	5021 => std_logic_vector(to_unsigned(42, 8)),
	5022 => std_logic_vector(to_unsigned(42, 8)),
	5023 => std_logic_vector(to_unsigned(42, 8)),
	5024 => std_logic_vector(to_unsigned(41, 8)),
	5025 => std_logic_vector(to_unsigned(41, 8)),
	5026 => std_logic_vector(to_unsigned(41, 8)),
	5027 => std_logic_vector(to_unsigned(41, 8)),
	5028 => std_logic_vector(to_unsigned(41, 8)),
	5029 => std_logic_vector(to_unsigned(41, 8)),
	5030 => std_logic_vector(to_unsigned(42, 8)),
	5031 => std_logic_vector(to_unsigned(42, 8)),
	5032 => std_logic_vector(to_unsigned(42, 8)),
	5033 => std_logic_vector(to_unsigned(41, 8)),
	5034 => std_logic_vector(to_unsigned(41, 8)),
	5035 => std_logic_vector(to_unsigned(41, 8)),
	5036 => std_logic_vector(to_unsigned(42, 8)),
	5037 => std_logic_vector(to_unsigned(41, 8)),
	5038 => std_logic_vector(to_unsigned(42, 8)),
	5039 => std_logic_vector(to_unsigned(42, 8)),
	5040 => std_logic_vector(to_unsigned(42, 8)),
	5041 => std_logic_vector(to_unsigned(41, 8)),
	5042 => std_logic_vector(to_unsigned(42, 8)),
	5043 => std_logic_vector(to_unsigned(41, 8)),
	5044 => std_logic_vector(to_unsigned(41, 8)),
	5045 => std_logic_vector(to_unsigned(41, 8)),
	5046 => std_logic_vector(to_unsigned(42, 8)),
	5047 => std_logic_vector(to_unsigned(42, 8)),
	5048 => std_logic_vector(to_unsigned(42, 8)),
	5049 => std_logic_vector(to_unsigned(42, 8)),
	5050 => std_logic_vector(to_unsigned(42, 8)),
	5051 => std_logic_vector(to_unsigned(41, 8)),
	5052 => std_logic_vector(to_unsigned(42, 8)),
	5053 => std_logic_vector(to_unsigned(41, 8)),
	5054 => std_logic_vector(to_unsigned(41, 8)),
	5055 => std_logic_vector(to_unsigned(41, 8)),
	5056 => std_logic_vector(to_unsigned(41, 8)),
	5057 => std_logic_vector(to_unsigned(41, 8)),
	5058 => std_logic_vector(to_unsigned(41, 8)),
	5059 => std_logic_vector(to_unsigned(42, 8)),
	5060 => std_logic_vector(to_unsigned(42, 8)),
	5061 => std_logic_vector(to_unsigned(42, 8)),
	5062 => std_logic_vector(to_unsigned(42, 8)),
	5063 => std_logic_vector(to_unsigned(42, 8)),
	5064 => std_logic_vector(to_unsigned(42, 8)),
	5065 => std_logic_vector(to_unsigned(41, 8)),
	5066 => std_logic_vector(to_unsigned(41, 8)),
	5067 => std_logic_vector(to_unsigned(41, 8)),
	5068 => std_logic_vector(to_unsigned(42, 8)),
	5069 => std_logic_vector(to_unsigned(41, 8)),
	5070 => std_logic_vector(to_unsigned(42, 8)),
	5071 => std_logic_vector(to_unsigned(42, 8)),
	5072 => std_logic_vector(to_unsigned(41, 8)),
	5073 => std_logic_vector(to_unsigned(41, 8)),
	5074 => std_logic_vector(to_unsigned(41, 8)),
	5075 => std_logic_vector(to_unsigned(41, 8)),
	5076 => std_logic_vector(to_unsigned(41, 8)),
	5077 => std_logic_vector(to_unsigned(42, 8)),
	5078 => std_logic_vector(to_unsigned(42, 8)),
	5079 => std_logic_vector(to_unsigned(42, 8)),
	5080 => std_logic_vector(to_unsigned(41, 8)),
	5081 => std_logic_vector(to_unsigned(42, 8)),
	5082 => std_logic_vector(to_unsigned(41, 8)),
	5083 => std_logic_vector(to_unsigned(41, 8)),
	5084 => std_logic_vector(to_unsigned(41, 8)),
	5085 => std_logic_vector(to_unsigned(41, 8)),
	5086 => std_logic_vector(to_unsigned(42, 8)),
	5087 => std_logic_vector(to_unsigned(41, 8)),
	5088 => std_logic_vector(to_unsigned(42, 8)),
	5089 => std_logic_vector(to_unsigned(42, 8)),
	5090 => std_logic_vector(to_unsigned(42, 8)),
	5091 => std_logic_vector(to_unsigned(42, 8)),
	5092 => std_logic_vector(to_unsigned(42, 8)),
	5093 => std_logic_vector(to_unsigned(41, 8)),
	5094 => std_logic_vector(to_unsigned(42, 8)),
	5095 => std_logic_vector(to_unsigned(42, 8)),
	5096 => std_logic_vector(to_unsigned(41, 8)),
	5097 => std_logic_vector(to_unsigned(42, 8)),
	5098 => std_logic_vector(to_unsigned(41, 8)),
	5099 => std_logic_vector(to_unsigned(42, 8)),
	5100 => std_logic_vector(to_unsigned(42, 8)),
	5101 => std_logic_vector(to_unsigned(41, 8)),
	5102 => std_logic_vector(to_unsigned(41, 8)),
	5103 => std_logic_vector(to_unsigned(42, 8)),
	5104 => std_logic_vector(to_unsigned(42, 8)),
	5105 => std_logic_vector(to_unsigned(41, 8)),
	5106 => std_logic_vector(to_unsigned(42, 8)),
	5107 => std_logic_vector(to_unsigned(41, 8)),
	5108 => std_logic_vector(to_unsigned(41, 8)),
	5109 => std_logic_vector(to_unsigned(41, 8)),
	5110 => std_logic_vector(to_unsigned(42, 8)),
	5111 => std_logic_vector(to_unsigned(41, 8)),
	5112 => std_logic_vector(to_unsigned(42, 8)),
	5113 => std_logic_vector(to_unsigned(42, 8)),
	5114 => std_logic_vector(to_unsigned(41, 8)),
	5115 => std_logic_vector(to_unsigned(41, 8)),
	5116 => std_logic_vector(to_unsigned(41, 8)),
	5117 => std_logic_vector(to_unsigned(42, 8)),
	5118 => std_logic_vector(to_unsigned(41, 8)),
	5119 => std_logic_vector(to_unsigned(42, 8)),
	5120 => std_logic_vector(to_unsigned(42, 8)),
	5121 => std_logic_vector(to_unsigned(42, 8)),
	5122 => std_logic_vector(to_unsigned(41, 8)),
	5123 => std_logic_vector(to_unsigned(41, 8)),
	5124 => std_logic_vector(to_unsigned(42, 8)),
	5125 => std_logic_vector(to_unsigned(42, 8)),
	5126 => std_logic_vector(to_unsigned(41, 8)),
	5127 => std_logic_vector(to_unsigned(41, 8)),
	5128 => std_logic_vector(to_unsigned(41, 8)),
	5129 => std_logic_vector(to_unsigned(41, 8)),
	5130 => std_logic_vector(to_unsigned(42, 8)),
	5131 => std_logic_vector(to_unsigned(41, 8)),
	5132 => std_logic_vector(to_unsigned(42, 8)),
	5133 => std_logic_vector(to_unsigned(42, 8)),
	5134 => std_logic_vector(to_unsigned(42, 8)),
	5135 => std_logic_vector(to_unsigned(41, 8)),
	5136 => std_logic_vector(to_unsigned(41, 8)),
	5137 => std_logic_vector(to_unsigned(42, 8)),
	5138 => std_logic_vector(to_unsigned(41, 8)),
	5139 => std_logic_vector(to_unsigned(42, 8)),
	5140 => std_logic_vector(to_unsigned(42, 8)),
	5141 => std_logic_vector(to_unsigned(41, 8)),
	5142 => std_logic_vector(to_unsigned(42, 8)),
	5143 => std_logic_vector(to_unsigned(41, 8)),
	5144 => std_logic_vector(to_unsigned(42, 8)),
	5145 => std_logic_vector(to_unsigned(42, 8)),
	5146 => std_logic_vector(to_unsigned(42, 8)),
	5147 => std_logic_vector(to_unsigned(41, 8)),
	5148 => std_logic_vector(to_unsigned(41, 8)),
	5149 => std_logic_vector(to_unsigned(42, 8)),
	5150 => std_logic_vector(to_unsigned(42, 8)),
	5151 => std_logic_vector(to_unsigned(41, 8)),
	5152 => std_logic_vector(to_unsigned(41, 8)),
	5153 => std_logic_vector(to_unsigned(41, 8)),
	5154 => std_logic_vector(to_unsigned(42, 8)),
	5155 => std_logic_vector(to_unsigned(42, 8)),
	5156 => std_logic_vector(to_unsigned(41, 8)),
	5157 => std_logic_vector(to_unsigned(41, 8)),
	5158 => std_logic_vector(to_unsigned(42, 8)),
	5159 => std_logic_vector(to_unsigned(41, 8)),
	5160 => std_logic_vector(to_unsigned(41, 8)),
	5161 => std_logic_vector(to_unsigned(42, 8)),
	5162 => std_logic_vector(to_unsigned(41, 8)),
	5163 => std_logic_vector(to_unsigned(41, 8)),
	5164 => std_logic_vector(to_unsigned(42, 8)),
	5165 => std_logic_vector(to_unsigned(42, 8)),
	5166 => std_logic_vector(to_unsigned(41, 8)),
	5167 => std_logic_vector(to_unsigned(42, 8)),
	5168 => std_logic_vector(to_unsigned(41, 8)),
	5169 => std_logic_vector(to_unsigned(41, 8)),
	5170 => std_logic_vector(to_unsigned(42, 8)),
	5171 => std_logic_vector(to_unsigned(41, 8)),
	5172 => std_logic_vector(to_unsigned(42, 8)),
	5173 => std_logic_vector(to_unsigned(41, 8)),
	5174 => std_logic_vector(to_unsigned(42, 8)),
	5175 => std_logic_vector(to_unsigned(42, 8)),
	5176 => std_logic_vector(to_unsigned(42, 8)),
	5177 => std_logic_vector(to_unsigned(41, 8)),
	5178 => std_logic_vector(to_unsigned(41, 8)),
	5179 => std_logic_vector(to_unsigned(41, 8)),
	5180 => std_logic_vector(to_unsigned(42, 8)),
	5181 => std_logic_vector(to_unsigned(41, 8)),
	5182 => std_logic_vector(to_unsigned(42, 8)),
	5183 => std_logic_vector(to_unsigned(41, 8)),
	5184 => std_logic_vector(to_unsigned(42, 8)),
	5185 => std_logic_vector(to_unsigned(41, 8)),
	5186 => std_logic_vector(to_unsigned(42, 8)),
	5187 => std_logic_vector(to_unsigned(42, 8)),
	5188 => std_logic_vector(to_unsigned(42, 8)),
	5189 => std_logic_vector(to_unsigned(41, 8)),
	5190 => std_logic_vector(to_unsigned(42, 8)),
	5191 => std_logic_vector(to_unsigned(41, 8)),
	5192 => std_logic_vector(to_unsigned(42, 8)),
	5193 => std_logic_vector(to_unsigned(42, 8)),
	5194 => std_logic_vector(to_unsigned(42, 8)),
	5195 => std_logic_vector(to_unsigned(42, 8)),
	5196 => std_logic_vector(to_unsigned(42, 8)),
	5197 => std_logic_vector(to_unsigned(41, 8)),
	5198 => std_logic_vector(to_unsigned(42, 8)),
	5199 => std_logic_vector(to_unsigned(42, 8)),
	5200 => std_logic_vector(to_unsigned(41, 8)),
	5201 => std_logic_vector(to_unsigned(42, 8)),
	5202 => std_logic_vector(to_unsigned(42, 8)),
	5203 => std_logic_vector(to_unsigned(41, 8)),
	5204 => std_logic_vector(to_unsigned(42, 8)),
	5205 => std_logic_vector(to_unsigned(41, 8)),
	5206 => std_logic_vector(to_unsigned(42, 8)),
	5207 => std_logic_vector(to_unsigned(42, 8)),
	5208 => std_logic_vector(to_unsigned(41, 8)),
	5209 => std_logic_vector(to_unsigned(42, 8)),
	5210 => std_logic_vector(to_unsigned(42, 8)),
	5211 => std_logic_vector(to_unsigned(42, 8)),
	5212 => std_logic_vector(to_unsigned(42, 8)),
	5213 => std_logic_vector(to_unsigned(41, 8)),
	5214 => std_logic_vector(to_unsigned(42, 8)),
	5215 => std_logic_vector(to_unsigned(41, 8)),
	5216 => std_logic_vector(to_unsigned(41, 8)),
	5217 => std_logic_vector(to_unsigned(41, 8)),
	5218 => std_logic_vector(to_unsigned(42, 8)),
	5219 => std_logic_vector(to_unsigned(42, 8)),
	5220 => std_logic_vector(to_unsigned(42, 8)),
	5221 => std_logic_vector(to_unsigned(42, 8)),
	5222 => std_logic_vector(to_unsigned(42, 8)),
	5223 => std_logic_vector(to_unsigned(41, 8)),
	5224 => std_logic_vector(to_unsigned(42, 8)),
	5225 => std_logic_vector(to_unsigned(42, 8)),
	5226 => std_logic_vector(to_unsigned(42, 8)),
	5227 => std_logic_vector(to_unsigned(41, 8)),
	5228 => std_logic_vector(to_unsigned(41, 8)),
	5229 => std_logic_vector(to_unsigned(42, 8)),
	5230 => std_logic_vector(to_unsigned(42, 8)),
	5231 => std_logic_vector(to_unsigned(41, 8)),
	5232 => std_logic_vector(to_unsigned(42, 8)),
	5233 => std_logic_vector(to_unsigned(42, 8)),
	5234 => std_logic_vector(to_unsigned(41, 8)),
	5235 => std_logic_vector(to_unsigned(42, 8)),
	5236 => std_logic_vector(to_unsigned(41, 8)),
	5237 => std_logic_vector(to_unsigned(41, 8)),
	5238 => std_logic_vector(to_unsigned(42, 8)),
	5239 => std_logic_vector(to_unsigned(42, 8)),
	5240 => std_logic_vector(to_unsigned(42, 8)),
	5241 => std_logic_vector(to_unsigned(41, 8)),
	5242 => std_logic_vector(to_unsigned(41, 8)),
	5243 => std_logic_vector(to_unsigned(41, 8)),
	5244 => std_logic_vector(to_unsigned(41, 8)),
	5245 => std_logic_vector(to_unsigned(42, 8)),
	5246 => std_logic_vector(to_unsigned(41, 8)),
	5247 => std_logic_vector(to_unsigned(41, 8)),
	5248 => std_logic_vector(to_unsigned(42, 8)),
	5249 => std_logic_vector(to_unsigned(42, 8)),
	5250 => std_logic_vector(to_unsigned(41, 8)),
	5251 => std_logic_vector(to_unsigned(41, 8)),
	5252 => std_logic_vector(to_unsigned(41, 8)),
	5253 => std_logic_vector(to_unsigned(41, 8)),
	5254 => std_logic_vector(to_unsigned(42, 8)),
	5255 => std_logic_vector(to_unsigned(42, 8)),
	5256 => std_logic_vector(to_unsigned(41, 8)),
	5257 => std_logic_vector(to_unsigned(42, 8)),
	5258 => std_logic_vector(to_unsigned(41, 8)),
	5259 => std_logic_vector(to_unsigned(41, 8)),
	5260 => std_logic_vector(to_unsigned(42, 8)),
	5261 => std_logic_vector(to_unsigned(42, 8)),
	5262 => std_logic_vector(to_unsigned(42, 8)),
	5263 => std_logic_vector(to_unsigned(42, 8)),
	5264 => std_logic_vector(to_unsigned(41, 8)),
	5265 => std_logic_vector(to_unsigned(42, 8)),
	5266 => std_logic_vector(to_unsigned(42, 8)),
	5267 => std_logic_vector(to_unsigned(42, 8)),
	5268 => std_logic_vector(to_unsigned(42, 8)),
	5269 => std_logic_vector(to_unsigned(41, 8)),
	5270 => std_logic_vector(to_unsigned(41, 8)),
	5271 => std_logic_vector(to_unsigned(41, 8)),
	5272 => std_logic_vector(to_unsigned(41, 8)),
	5273 => std_logic_vector(to_unsigned(41, 8)),
	5274 => std_logic_vector(to_unsigned(42, 8)),
	5275 => std_logic_vector(to_unsigned(41, 8)),
	5276 => std_logic_vector(to_unsigned(42, 8)),
	5277 => std_logic_vector(to_unsigned(41, 8)),
	5278 => std_logic_vector(to_unsigned(41, 8)),
	5279 => std_logic_vector(to_unsigned(41, 8)),
	5280 => std_logic_vector(to_unsigned(41, 8)),
	5281 => std_logic_vector(to_unsigned(42, 8)),
	5282 => std_logic_vector(to_unsigned(42, 8)),
	5283 => std_logic_vector(to_unsigned(41, 8)),
	5284 => std_logic_vector(to_unsigned(42, 8)),
	5285 => std_logic_vector(to_unsigned(41, 8)),
	5286 => std_logic_vector(to_unsigned(41, 8)),
	5287 => std_logic_vector(to_unsigned(41, 8)),
	5288 => std_logic_vector(to_unsigned(41, 8)),
	5289 => std_logic_vector(to_unsigned(42, 8)),
	5290 => std_logic_vector(to_unsigned(42, 8)),
	5291 => std_logic_vector(to_unsigned(41, 8)),
	5292 => std_logic_vector(to_unsigned(41, 8)),
	5293 => std_logic_vector(to_unsigned(41, 8)),
	5294 => std_logic_vector(to_unsigned(42, 8)),
	5295 => std_logic_vector(to_unsigned(42, 8)),
	5296 => std_logic_vector(to_unsigned(42, 8)),
	5297 => std_logic_vector(to_unsigned(42, 8)),
	5298 => std_logic_vector(to_unsigned(41, 8)),
	5299 => std_logic_vector(to_unsigned(42, 8)),
	5300 => std_logic_vector(to_unsigned(41, 8)),
	5301 => std_logic_vector(to_unsigned(41, 8)),
	5302 => std_logic_vector(to_unsigned(42, 8)),
	5303 => std_logic_vector(to_unsigned(41, 8)),
	5304 => std_logic_vector(to_unsigned(42, 8)),
	5305 => std_logic_vector(to_unsigned(41, 8)),
	5306 => std_logic_vector(to_unsigned(42, 8)),
	5307 => std_logic_vector(to_unsigned(41, 8)),
	5308 => std_logic_vector(to_unsigned(41, 8)),
	5309 => std_logic_vector(to_unsigned(41, 8)),
	5310 => std_logic_vector(to_unsigned(42, 8)),
	5311 => std_logic_vector(to_unsigned(41, 8)),
	5312 => std_logic_vector(to_unsigned(41, 8)),
	5313 => std_logic_vector(to_unsigned(42, 8)),
	5314 => std_logic_vector(to_unsigned(41, 8)),
	5315 => std_logic_vector(to_unsigned(41, 8)),
	5316 => std_logic_vector(to_unsigned(41, 8)),
	5317 => std_logic_vector(to_unsigned(41, 8)),
	5318 => std_logic_vector(to_unsigned(41, 8)),
	5319 => std_logic_vector(to_unsigned(42, 8)),
	5320 => std_logic_vector(to_unsigned(42, 8)),
	5321 => std_logic_vector(to_unsigned(42, 8)),
	5322 => std_logic_vector(to_unsigned(41, 8)),
	5323 => std_logic_vector(to_unsigned(42, 8)),
	5324 => std_logic_vector(to_unsigned(42, 8)),
	5325 => std_logic_vector(to_unsigned(41, 8)),
	5326 => std_logic_vector(to_unsigned(41, 8)),
	5327 => std_logic_vector(to_unsigned(41, 8)),
	5328 => std_logic_vector(to_unsigned(41, 8)),
	5329 => std_logic_vector(to_unsigned(41, 8)),
	5330 => std_logic_vector(to_unsigned(41, 8)),
	5331 => std_logic_vector(to_unsigned(41, 8)),
	5332 => std_logic_vector(to_unsigned(42, 8)),
	5333 => std_logic_vector(to_unsigned(42, 8)),
	5334 => std_logic_vector(to_unsigned(41, 8)),
	5335 => std_logic_vector(to_unsigned(41, 8)),
	5336 => std_logic_vector(to_unsigned(41, 8)),
	5337 => std_logic_vector(to_unsigned(42, 8)),
	5338 => std_logic_vector(to_unsigned(41, 8)),
	5339 => std_logic_vector(to_unsigned(41, 8)),
	5340 => std_logic_vector(to_unsigned(42, 8)),
	5341 => std_logic_vector(to_unsigned(42, 8)),
	5342 => std_logic_vector(to_unsigned(42, 8)),
	5343 => std_logic_vector(to_unsigned(42, 8)),
	5344 => std_logic_vector(to_unsigned(42, 8)),
	5345 => std_logic_vector(to_unsigned(41, 8)),
	5346 => std_logic_vector(to_unsigned(41, 8)),
	5347 => std_logic_vector(to_unsigned(41, 8)),
	5348 => std_logic_vector(to_unsigned(41, 8)),
	5349 => std_logic_vector(to_unsigned(42, 8)),
	5350 => std_logic_vector(to_unsigned(42, 8)),
	5351 => std_logic_vector(to_unsigned(42, 8)),
	5352 => std_logic_vector(to_unsigned(41, 8)),
	5353 => std_logic_vector(to_unsigned(41, 8)),
	5354 => std_logic_vector(to_unsigned(42, 8)),
	5355 => std_logic_vector(to_unsigned(42, 8)),
	5356 => std_logic_vector(to_unsigned(41, 8)),
	5357 => std_logic_vector(to_unsigned(41, 8)),
	5358 => std_logic_vector(to_unsigned(41, 8)),
	5359 => std_logic_vector(to_unsigned(41, 8)),
	5360 => std_logic_vector(to_unsigned(42, 8)),
	5361 => std_logic_vector(to_unsigned(42, 8)),
	5362 => std_logic_vector(to_unsigned(42, 8)),
	5363 => std_logic_vector(to_unsigned(41, 8)),
	5364 => std_logic_vector(to_unsigned(41, 8)),
	5365 => std_logic_vector(to_unsigned(42, 8)),
	5366 => std_logic_vector(to_unsigned(41, 8)),
	5367 => std_logic_vector(to_unsigned(41, 8)),
	5368 => std_logic_vector(to_unsigned(41, 8)),
	5369 => std_logic_vector(to_unsigned(41, 8)),
	5370 => std_logic_vector(to_unsigned(41, 8)),
	5371 => std_logic_vector(to_unsigned(42, 8)),
	5372 => std_logic_vector(to_unsigned(41, 8)),
	5373 => std_logic_vector(to_unsigned(41, 8)),
	5374 => std_logic_vector(to_unsigned(42, 8)),
	5375 => std_logic_vector(to_unsigned(41, 8)),
	5376 => std_logic_vector(to_unsigned(41, 8)),
	5377 => std_logic_vector(to_unsigned(41, 8)),
	5378 => std_logic_vector(to_unsigned(42, 8)),
	5379 => std_logic_vector(to_unsigned(42, 8)),
	5380 => std_logic_vector(to_unsigned(41, 8)),
	5381 => std_logic_vector(to_unsigned(42, 8)),
	5382 => std_logic_vector(to_unsigned(41, 8)),
	5383 => std_logic_vector(to_unsigned(42, 8)),
	5384 => std_logic_vector(to_unsigned(42, 8)),
	5385 => std_logic_vector(to_unsigned(41, 8)),
	5386 => std_logic_vector(to_unsigned(42, 8)),
	5387 => std_logic_vector(to_unsigned(42, 8)),
	5388 => std_logic_vector(to_unsigned(41, 8)),
	5389 => std_logic_vector(to_unsigned(42, 8)),
	5390 => std_logic_vector(to_unsigned(42, 8)),
	5391 => std_logic_vector(to_unsigned(42, 8)),
	5392 => std_logic_vector(to_unsigned(41, 8)),
	5393 => std_logic_vector(to_unsigned(41, 8)),
	5394 => std_logic_vector(to_unsigned(41, 8)),
	5395 => std_logic_vector(to_unsigned(41, 8)),
	5396 => std_logic_vector(to_unsigned(42, 8)),
	5397 => std_logic_vector(to_unsigned(42, 8)),
	5398 => std_logic_vector(to_unsigned(41, 8)),
	5399 => std_logic_vector(to_unsigned(41, 8)),
	5400 => std_logic_vector(to_unsigned(41, 8)),
	5401 => std_logic_vector(to_unsigned(42, 8)),
	5402 => std_logic_vector(to_unsigned(42, 8)),
	5403 => std_logic_vector(to_unsigned(41, 8)),
	5404 => std_logic_vector(to_unsigned(41, 8)),
	5405 => std_logic_vector(to_unsigned(42, 8)),
	5406 => std_logic_vector(to_unsigned(41, 8)),
	5407 => std_logic_vector(to_unsigned(42, 8)),
	5408 => std_logic_vector(to_unsigned(41, 8)),
	5409 => std_logic_vector(to_unsigned(42, 8)),
	5410 => std_logic_vector(to_unsigned(42, 8)),
	5411 => std_logic_vector(to_unsigned(41, 8)),
	5412 => std_logic_vector(to_unsigned(41, 8)),
	5413 => std_logic_vector(to_unsigned(41, 8)),
	5414 => std_logic_vector(to_unsigned(41, 8)),
	5415 => std_logic_vector(to_unsigned(41, 8)),
	5416 => std_logic_vector(to_unsigned(41, 8)),
	5417 => std_logic_vector(to_unsigned(41, 8)),
	5418 => std_logic_vector(to_unsigned(41, 8)),
	5419 => std_logic_vector(to_unsigned(42, 8)),
	5420 => std_logic_vector(to_unsigned(42, 8)),
	5421 => std_logic_vector(to_unsigned(42, 8)),
	5422 => std_logic_vector(to_unsigned(41, 8)),
	5423 => std_logic_vector(to_unsigned(41, 8)),
	5424 => std_logic_vector(to_unsigned(41, 8)),
	5425 => std_logic_vector(to_unsigned(42, 8)),
	5426 => std_logic_vector(to_unsigned(42, 8)),
	5427 => std_logic_vector(to_unsigned(42, 8)),
	5428 => std_logic_vector(to_unsigned(42, 8)),
	5429 => std_logic_vector(to_unsigned(41, 8)),
	5430 => std_logic_vector(to_unsigned(41, 8)),
	5431 => std_logic_vector(to_unsigned(41, 8)),
	5432 => std_logic_vector(to_unsigned(41, 8)),
	5433 => std_logic_vector(to_unsigned(41, 8)),
	5434 => std_logic_vector(to_unsigned(41, 8)),
	5435 => std_logic_vector(to_unsigned(41, 8)),
	5436 => std_logic_vector(to_unsigned(42, 8)),
	5437 => std_logic_vector(to_unsigned(41, 8)),
	5438 => std_logic_vector(to_unsigned(42, 8)),
	5439 => std_logic_vector(to_unsigned(42, 8)),
	5440 => std_logic_vector(to_unsigned(42, 8)),
	5441 => std_logic_vector(to_unsigned(42, 8)),
	5442 => std_logic_vector(to_unsigned(41, 8)),
	5443 => std_logic_vector(to_unsigned(42, 8)),
	5444 => std_logic_vector(to_unsigned(42, 8)),
	5445 => std_logic_vector(to_unsigned(41, 8)),
	5446 => std_logic_vector(to_unsigned(41, 8)),
	5447 => std_logic_vector(to_unsigned(41, 8)),
	5448 => std_logic_vector(to_unsigned(41, 8)),
	5449 => std_logic_vector(to_unsigned(41, 8)),
	5450 => std_logic_vector(to_unsigned(42, 8)),
	5451 => std_logic_vector(to_unsigned(41, 8)),
	5452 => std_logic_vector(to_unsigned(42, 8)),
	5453 => std_logic_vector(to_unsigned(41, 8)),
	5454 => std_logic_vector(to_unsigned(42, 8)),
	5455 => std_logic_vector(to_unsigned(41, 8)),
	5456 => std_logic_vector(to_unsigned(41, 8)),
	5457 => std_logic_vector(to_unsigned(42, 8)),
	5458 => std_logic_vector(to_unsigned(42, 8)),
	5459 => std_logic_vector(to_unsigned(42, 8)),
	5460 => std_logic_vector(to_unsigned(41, 8)),
	5461 => std_logic_vector(to_unsigned(42, 8)),
	5462 => std_logic_vector(to_unsigned(42, 8)),
	5463 => std_logic_vector(to_unsigned(42, 8)),
	5464 => std_logic_vector(to_unsigned(42, 8)),
	5465 => std_logic_vector(to_unsigned(42, 8)),
	5466 => std_logic_vector(to_unsigned(41, 8)),
	5467 => std_logic_vector(to_unsigned(42, 8)),
	5468 => std_logic_vector(to_unsigned(42, 8)),
	5469 => std_logic_vector(to_unsigned(41, 8)),
	5470 => std_logic_vector(to_unsigned(41, 8)),
	5471 => std_logic_vector(to_unsigned(42, 8)),
	5472 => std_logic_vector(to_unsigned(42, 8)),
	5473 => std_logic_vector(to_unsigned(41, 8)),
	5474 => std_logic_vector(to_unsigned(42, 8)),
	5475 => std_logic_vector(to_unsigned(42, 8)),
	5476 => std_logic_vector(to_unsigned(42, 8)),
	5477 => std_logic_vector(to_unsigned(42, 8)),
	5478 => std_logic_vector(to_unsigned(42, 8)),
	5479 => std_logic_vector(to_unsigned(42, 8)),
	5480 => std_logic_vector(to_unsigned(42, 8)),
	5481 => std_logic_vector(to_unsigned(41, 8)),
	5482 => std_logic_vector(to_unsigned(41, 8)),
	5483 => std_logic_vector(to_unsigned(41, 8)),
	5484 => std_logic_vector(to_unsigned(42, 8)),
	5485 => std_logic_vector(to_unsigned(42, 8)),
	5486 => std_logic_vector(to_unsigned(42, 8)),
	5487 => std_logic_vector(to_unsigned(41, 8)),
	5488 => std_logic_vector(to_unsigned(42, 8)),
	5489 => std_logic_vector(to_unsigned(41, 8)),
	5490 => std_logic_vector(to_unsigned(42, 8)),
	5491 => std_logic_vector(to_unsigned(42, 8)),
	5492 => std_logic_vector(to_unsigned(42, 8)),
	5493 => std_logic_vector(to_unsigned(42, 8)),
	5494 => std_logic_vector(to_unsigned(41, 8)),
	5495 => std_logic_vector(to_unsigned(42, 8)),
	5496 => std_logic_vector(to_unsigned(41, 8)),
	5497 => std_logic_vector(to_unsigned(42, 8)),
	5498 => std_logic_vector(to_unsigned(41, 8)),
	5499 => std_logic_vector(to_unsigned(42, 8)),
	5500 => std_logic_vector(to_unsigned(41, 8)),
	5501 => std_logic_vector(to_unsigned(41, 8)),
	5502 => std_logic_vector(to_unsigned(42, 8)),
	5503 => std_logic_vector(to_unsigned(42, 8)),
	5504 => std_logic_vector(to_unsigned(41, 8)),
	5505 => std_logic_vector(to_unsigned(42, 8)),
	5506 => std_logic_vector(to_unsigned(41, 8)),
	5507 => std_logic_vector(to_unsigned(42, 8)),
	5508 => std_logic_vector(to_unsigned(41, 8)),
	5509 => std_logic_vector(to_unsigned(41, 8)),
	5510 => std_logic_vector(to_unsigned(42, 8)),
	5511 => std_logic_vector(to_unsigned(42, 8)),
	5512 => std_logic_vector(to_unsigned(41, 8)),
	5513 => std_logic_vector(to_unsigned(42, 8)),
	5514 => std_logic_vector(to_unsigned(42, 8)),
	5515 => std_logic_vector(to_unsigned(41, 8)),
	5516 => std_logic_vector(to_unsigned(41, 8)),
	5517 => std_logic_vector(to_unsigned(41, 8)),
	5518 => std_logic_vector(to_unsigned(41, 8)),
	5519 => std_logic_vector(to_unsigned(42, 8)),
	5520 => std_logic_vector(to_unsigned(42, 8)),
	5521 => std_logic_vector(to_unsigned(41, 8)),
	5522 => std_logic_vector(to_unsigned(42, 8)),
	5523 => std_logic_vector(to_unsigned(41, 8)),
	5524 => std_logic_vector(to_unsigned(41, 8)),
	5525 => std_logic_vector(to_unsigned(42, 8)),
	5526 => std_logic_vector(to_unsigned(42, 8)),
	5527 => std_logic_vector(to_unsigned(41, 8)),
	5528 => std_logic_vector(to_unsigned(41, 8)),
	5529 => std_logic_vector(to_unsigned(41, 8)),
	5530 => std_logic_vector(to_unsigned(41, 8)),
	5531 => std_logic_vector(to_unsigned(42, 8)),
	5532 => std_logic_vector(to_unsigned(42, 8)),
	5533 => std_logic_vector(to_unsigned(41, 8)),
	5534 => std_logic_vector(to_unsigned(41, 8)),
	5535 => std_logic_vector(to_unsigned(42, 8)),
	5536 => std_logic_vector(to_unsigned(41, 8)),
	5537 => std_logic_vector(to_unsigned(41, 8)),
	5538 => std_logic_vector(to_unsigned(41, 8)),
	5539 => std_logic_vector(to_unsigned(42, 8)),
	5540 => std_logic_vector(to_unsigned(42, 8)),
	5541 => std_logic_vector(to_unsigned(42, 8)),
	5542 => std_logic_vector(to_unsigned(41, 8)),
	5543 => std_logic_vector(to_unsigned(41, 8)),
	5544 => std_logic_vector(to_unsigned(42, 8)),
	5545 => std_logic_vector(to_unsigned(41, 8)),
	5546 => std_logic_vector(to_unsigned(42, 8)),
	5547 => std_logic_vector(to_unsigned(42, 8)),
	5548 => std_logic_vector(to_unsigned(42, 8)),
	5549 => std_logic_vector(to_unsigned(41, 8)),
	5550 => std_logic_vector(to_unsigned(41, 8)),
	5551 => std_logic_vector(to_unsigned(41, 8)),
	5552 => std_logic_vector(to_unsigned(41, 8)),
	5553 => std_logic_vector(to_unsigned(42, 8)),
	5554 => std_logic_vector(to_unsigned(42, 8)),
	5555 => std_logic_vector(to_unsigned(41, 8)),
	5556 => std_logic_vector(to_unsigned(42, 8)),
	5557 => std_logic_vector(to_unsigned(42, 8)),
	5558 => std_logic_vector(to_unsigned(42, 8)),
	5559 => std_logic_vector(to_unsigned(41, 8)),
	5560 => std_logic_vector(to_unsigned(41, 8)),
	5561 => std_logic_vector(to_unsigned(42, 8)),
	5562 => std_logic_vector(to_unsigned(41, 8)),
	5563 => std_logic_vector(to_unsigned(41, 8)),
	5564 => std_logic_vector(to_unsigned(41, 8)),
	5565 => std_logic_vector(to_unsigned(41, 8)),
	5566 => std_logic_vector(to_unsigned(41, 8)),
	5567 => std_logic_vector(to_unsigned(42, 8)),
	5568 => std_logic_vector(to_unsigned(41, 8)),
	5569 => std_logic_vector(to_unsigned(42, 8)),
	5570 => std_logic_vector(to_unsigned(42, 8)),
	5571 => std_logic_vector(to_unsigned(42, 8)),
	5572 => std_logic_vector(to_unsigned(42, 8)),
	5573 => std_logic_vector(to_unsigned(42, 8)),
	5574 => std_logic_vector(to_unsigned(41, 8)),
	5575 => std_logic_vector(to_unsigned(41, 8)),
	5576 => std_logic_vector(to_unsigned(41, 8)),
	5577 => std_logic_vector(to_unsigned(42, 8)),
	5578 => std_logic_vector(to_unsigned(41, 8)),
	5579 => std_logic_vector(to_unsigned(41, 8)),
	5580 => std_logic_vector(to_unsigned(42, 8)),
	5581 => std_logic_vector(to_unsigned(42, 8)),
	5582 => std_logic_vector(to_unsigned(42, 8)),
	5583 => std_logic_vector(to_unsigned(41, 8)),
	5584 => std_logic_vector(to_unsigned(42, 8)),
	5585 => std_logic_vector(to_unsigned(42, 8)),
	5586 => std_logic_vector(to_unsigned(41, 8)),
	5587 => std_logic_vector(to_unsigned(41, 8)),
	5588 => std_logic_vector(to_unsigned(41, 8)),
	5589 => std_logic_vector(to_unsigned(41, 8)),
	5590 => std_logic_vector(to_unsigned(42, 8)),
	5591 => std_logic_vector(to_unsigned(41, 8)),
	5592 => std_logic_vector(to_unsigned(41, 8)),
	5593 => std_logic_vector(to_unsigned(42, 8)),
	5594 => std_logic_vector(to_unsigned(42, 8)),
	5595 => std_logic_vector(to_unsigned(42, 8)),
	5596 => std_logic_vector(to_unsigned(41, 8)),
	5597 => std_logic_vector(to_unsigned(42, 8)),
	5598 => std_logic_vector(to_unsigned(41, 8)),
	5599 => std_logic_vector(to_unsigned(42, 8)),
	5600 => std_logic_vector(to_unsigned(41, 8)),
	5601 => std_logic_vector(to_unsigned(42, 8)),
	5602 => std_logic_vector(to_unsigned(41, 8)),
	5603 => std_logic_vector(to_unsigned(42, 8)),
	5604 => std_logic_vector(to_unsigned(41, 8)),
	5605 => std_logic_vector(to_unsigned(42, 8)),
	5606 => std_logic_vector(to_unsigned(41, 8)),
	5607 => std_logic_vector(to_unsigned(42, 8)),
	5608 => std_logic_vector(to_unsigned(42, 8)),
	5609 => std_logic_vector(to_unsigned(42, 8)),
	5610 => std_logic_vector(to_unsigned(41, 8)),
	5611 => std_logic_vector(to_unsigned(41, 8)),
	5612 => std_logic_vector(to_unsigned(42, 8)),
	5613 => std_logic_vector(to_unsigned(41, 8)),
	5614 => std_logic_vector(to_unsigned(41, 8)),
	5615 => std_logic_vector(to_unsigned(41, 8)),
	5616 => std_logic_vector(to_unsigned(41, 8)),
	5617 => std_logic_vector(to_unsigned(41, 8)),
	5618 => std_logic_vector(to_unsigned(42, 8)),
	5619 => std_logic_vector(to_unsigned(41, 8)),
	5620 => std_logic_vector(to_unsigned(42, 8)),
	5621 => std_logic_vector(to_unsigned(41, 8)),
	5622 => std_logic_vector(to_unsigned(42, 8)),
	5623 => std_logic_vector(to_unsigned(42, 8)),
	5624 => std_logic_vector(to_unsigned(42, 8)),
	5625 => std_logic_vector(to_unsigned(42, 8)),
	5626 => std_logic_vector(to_unsigned(41, 8)),
	5627 => std_logic_vector(to_unsigned(42, 8)),
	5628 => std_logic_vector(to_unsigned(42, 8)),
	5629 => std_logic_vector(to_unsigned(41, 8)),
	5630 => std_logic_vector(to_unsigned(41, 8)),
	5631 => std_logic_vector(to_unsigned(41, 8)),
	5632 => std_logic_vector(to_unsigned(41, 8)),
	5633 => std_logic_vector(to_unsigned(42, 8)),
	5634 => std_logic_vector(to_unsigned(41, 8)),
	5635 => std_logic_vector(to_unsigned(41, 8)),
	5636 => std_logic_vector(to_unsigned(42, 8)),
	5637 => std_logic_vector(to_unsigned(41, 8)),
	5638 => std_logic_vector(to_unsigned(42, 8)),
	5639 => std_logic_vector(to_unsigned(41, 8)),
	5640 => std_logic_vector(to_unsigned(41, 8)),
	5641 => std_logic_vector(to_unsigned(42, 8)),
	5642 => std_logic_vector(to_unsigned(41, 8)),
	5643 => std_logic_vector(to_unsigned(41, 8)),
	5644 => std_logic_vector(to_unsigned(41, 8)),
	5645 => std_logic_vector(to_unsigned(41, 8)),
	5646 => std_logic_vector(to_unsigned(42, 8)),
	5647 => std_logic_vector(to_unsigned(42, 8)),
	5648 => std_logic_vector(to_unsigned(41, 8)),
	5649 => std_logic_vector(to_unsigned(41, 8)),
	5650 => std_logic_vector(to_unsigned(42, 8)),
	5651 => std_logic_vector(to_unsigned(42, 8)),
	5652 => std_logic_vector(to_unsigned(42, 8)),
	5653 => std_logic_vector(to_unsigned(41, 8)),
	5654 => std_logic_vector(to_unsigned(41, 8)),
	5655 => std_logic_vector(to_unsigned(41, 8)),
	5656 => std_logic_vector(to_unsigned(42, 8)),
	5657 => std_logic_vector(to_unsigned(41, 8)),
	5658 => std_logic_vector(to_unsigned(42, 8)),
	5659 => std_logic_vector(to_unsigned(41, 8)),
	5660 => std_logic_vector(to_unsigned(42, 8)),
	5661 => std_logic_vector(to_unsigned(41, 8)),
	5662 => std_logic_vector(to_unsigned(42, 8)),
	5663 => std_logic_vector(to_unsigned(42, 8)),
	5664 => std_logic_vector(to_unsigned(42, 8)),
	5665 => std_logic_vector(to_unsigned(42, 8)),
	5666 => std_logic_vector(to_unsigned(42, 8)),
	5667 => std_logic_vector(to_unsigned(42, 8)),
	5668 => std_logic_vector(to_unsigned(42, 8)),
	5669 => std_logic_vector(to_unsigned(42, 8)),
	5670 => std_logic_vector(to_unsigned(42, 8)),
	5671 => std_logic_vector(to_unsigned(42, 8)),
	5672 => std_logic_vector(to_unsigned(41, 8)),
	5673 => std_logic_vector(to_unsigned(41, 8)),
	5674 => std_logic_vector(to_unsigned(41, 8)),
	5675 => std_logic_vector(to_unsigned(42, 8)),
	5676 => std_logic_vector(to_unsigned(42, 8)),
	5677 => std_logic_vector(to_unsigned(41, 8)),
	5678 => std_logic_vector(to_unsigned(42, 8)),
	5679 => std_logic_vector(to_unsigned(41, 8)),
	5680 => std_logic_vector(to_unsigned(41, 8)),
	5681 => std_logic_vector(to_unsigned(42, 8)),
	5682 => std_logic_vector(to_unsigned(42, 8)),
	5683 => std_logic_vector(to_unsigned(42, 8)),
	5684 => std_logic_vector(to_unsigned(42, 8)),
	5685 => std_logic_vector(to_unsigned(42, 8)),
	5686 => std_logic_vector(to_unsigned(42, 8)),
	5687 => std_logic_vector(to_unsigned(41, 8)),
	5688 => std_logic_vector(to_unsigned(41, 8)),
	5689 => std_logic_vector(to_unsigned(41, 8)),
	5690 => std_logic_vector(to_unsigned(41, 8)),
	5691 => std_logic_vector(to_unsigned(42, 8)),
	5692 => std_logic_vector(to_unsigned(41, 8)),
	5693 => std_logic_vector(to_unsigned(42, 8)),
	5694 => std_logic_vector(to_unsigned(42, 8)),
	5695 => std_logic_vector(to_unsigned(41, 8)),
	5696 => std_logic_vector(to_unsigned(41, 8)),
	5697 => std_logic_vector(to_unsigned(41, 8)),
	5698 => std_logic_vector(to_unsigned(41, 8)),
	5699 => std_logic_vector(to_unsigned(41, 8)),
	5700 => std_logic_vector(to_unsigned(41, 8)),
	5701 => std_logic_vector(to_unsigned(41, 8)),
	5702 => std_logic_vector(to_unsigned(42, 8)),
	5703 => std_logic_vector(to_unsigned(41, 8)),
	5704 => std_logic_vector(to_unsigned(41, 8)),
	5705 => std_logic_vector(to_unsigned(41, 8)),
	5706 => std_logic_vector(to_unsigned(42, 8)),
	5707 => std_logic_vector(to_unsigned(41, 8)),
	5708 => std_logic_vector(to_unsigned(41, 8)),
	5709 => std_logic_vector(to_unsigned(42, 8)),
	5710 => std_logic_vector(to_unsigned(41, 8)),
	5711 => std_logic_vector(to_unsigned(41, 8)),
	5712 => std_logic_vector(to_unsigned(42, 8)),
	5713 => std_logic_vector(to_unsigned(42, 8)),
	5714 => std_logic_vector(to_unsigned(41, 8)),
	5715 => std_logic_vector(to_unsigned(41, 8)),
	5716 => std_logic_vector(to_unsigned(42, 8)),
	5717 => std_logic_vector(to_unsigned(41, 8)),
	5718 => std_logic_vector(to_unsigned(41, 8)),
	5719 => std_logic_vector(to_unsigned(42, 8)),
	5720 => std_logic_vector(to_unsigned(41, 8)),
	5721 => std_logic_vector(to_unsigned(42, 8)),
	5722 => std_logic_vector(to_unsigned(41, 8)),
	5723 => std_logic_vector(to_unsigned(41, 8)),
	5724 => std_logic_vector(to_unsigned(41, 8)),
	5725 => std_logic_vector(to_unsigned(42, 8)),
	5726 => std_logic_vector(to_unsigned(41, 8)),
	5727 => std_logic_vector(to_unsigned(42, 8)),
	5728 => std_logic_vector(to_unsigned(41, 8)),
	5729 => std_logic_vector(to_unsigned(41, 8)),
	5730 => std_logic_vector(to_unsigned(42, 8)),
	5731 => std_logic_vector(to_unsigned(42, 8)),
	5732 => std_logic_vector(to_unsigned(42, 8)),
	5733 => std_logic_vector(to_unsigned(42, 8)),
	5734 => std_logic_vector(to_unsigned(42, 8)),
	5735 => std_logic_vector(to_unsigned(41, 8)),
	5736 => std_logic_vector(to_unsigned(42, 8)),
	5737 => std_logic_vector(to_unsigned(42, 8)),
	5738 => std_logic_vector(to_unsigned(42, 8)),
	5739 => std_logic_vector(to_unsigned(41, 8)),
	5740 => std_logic_vector(to_unsigned(42, 8)),
	5741 => std_logic_vector(to_unsigned(42, 8)),
	5742 => std_logic_vector(to_unsigned(41, 8)),
	5743 => std_logic_vector(to_unsigned(42, 8)),
	5744 => std_logic_vector(to_unsigned(42, 8)),
	5745 => std_logic_vector(to_unsigned(41, 8)),
	5746 => std_logic_vector(to_unsigned(41, 8)),
	5747 => std_logic_vector(to_unsigned(42, 8)),
	5748 => std_logic_vector(to_unsigned(42, 8)),
	5749 => std_logic_vector(to_unsigned(41, 8)),
	5750 => std_logic_vector(to_unsigned(41, 8)),
	5751 => std_logic_vector(to_unsigned(41, 8)),
	5752 => std_logic_vector(to_unsigned(41, 8)),
	5753 => std_logic_vector(to_unsigned(41, 8)),
	5754 => std_logic_vector(to_unsigned(42, 8)),
	5755 => std_logic_vector(to_unsigned(42, 8)),
	5756 => std_logic_vector(to_unsigned(42, 8)),
	5757 => std_logic_vector(to_unsigned(41, 8)),
	5758 => std_logic_vector(to_unsigned(42, 8)),
	5759 => std_logic_vector(to_unsigned(42, 8)),
	5760 => std_logic_vector(to_unsigned(41, 8)),
	5761 => std_logic_vector(to_unsigned(42, 8)),
	5762 => std_logic_vector(to_unsigned(41, 8)),
	5763 => std_logic_vector(to_unsigned(42, 8)),
	5764 => std_logic_vector(to_unsigned(41, 8)),
	5765 => std_logic_vector(to_unsigned(41, 8)),
	5766 => std_logic_vector(to_unsigned(42, 8)),
	5767 => std_logic_vector(to_unsigned(42, 8)),
	5768 => std_logic_vector(to_unsigned(42, 8)),
	5769 => std_logic_vector(to_unsigned(42, 8)),
	5770 => std_logic_vector(to_unsigned(41, 8)),
	5771 => std_logic_vector(to_unsigned(41, 8)),
	5772 => std_logic_vector(to_unsigned(42, 8)),
	5773 => std_logic_vector(to_unsigned(41, 8)),
	5774 => std_logic_vector(to_unsigned(41, 8)),
	5775 => std_logic_vector(to_unsigned(41, 8)),
	5776 => std_logic_vector(to_unsigned(41, 8)),
	5777 => std_logic_vector(to_unsigned(41, 8)),
	5778 => std_logic_vector(to_unsigned(42, 8)),
	5779 => std_logic_vector(to_unsigned(41, 8)),
	5780 => std_logic_vector(to_unsigned(42, 8)),
	5781 => std_logic_vector(to_unsigned(41, 8)),
	5782 => std_logic_vector(to_unsigned(41, 8)),
	5783 => std_logic_vector(to_unsigned(41, 8)),
	5784 => std_logic_vector(to_unsigned(41, 8)),
	5785 => std_logic_vector(to_unsigned(42, 8)),
	5786 => std_logic_vector(to_unsigned(42, 8)),
	5787 => std_logic_vector(to_unsigned(41, 8)),
	5788 => std_logic_vector(to_unsigned(42, 8)),
	5789 => std_logic_vector(to_unsigned(41, 8)),
	5790 => std_logic_vector(to_unsigned(41, 8)),
	5791 => std_logic_vector(to_unsigned(41, 8)),
	5792 => std_logic_vector(to_unsigned(42, 8)),
	5793 => std_logic_vector(to_unsigned(41, 8)),
	5794 => std_logic_vector(to_unsigned(42, 8)),
	5795 => std_logic_vector(to_unsigned(41, 8)),
	5796 => std_logic_vector(to_unsigned(41, 8)),
	5797 => std_logic_vector(to_unsigned(42, 8)),
	5798 => std_logic_vector(to_unsigned(42, 8)),
	5799 => std_logic_vector(to_unsigned(41, 8)),
	5800 => std_logic_vector(to_unsigned(42, 8)),
	5801 => std_logic_vector(to_unsigned(41, 8)),
	5802 => std_logic_vector(to_unsigned(41, 8)),
	5803 => std_logic_vector(to_unsigned(41, 8)),
	5804 => std_logic_vector(to_unsigned(42, 8)),
	5805 => std_logic_vector(to_unsigned(42, 8)),
	5806 => std_logic_vector(to_unsigned(41, 8)),
	5807 => std_logic_vector(to_unsigned(42, 8)),
	5808 => std_logic_vector(to_unsigned(42, 8)),
	5809 => std_logic_vector(to_unsigned(41, 8)),
	5810 => std_logic_vector(to_unsigned(42, 8)),
	5811 => std_logic_vector(to_unsigned(42, 8)),
	5812 => std_logic_vector(to_unsigned(41, 8)),
	5813 => std_logic_vector(to_unsigned(41, 8)),
	5814 => std_logic_vector(to_unsigned(41, 8)),
	5815 => std_logic_vector(to_unsigned(41, 8)),
	5816 => std_logic_vector(to_unsigned(41, 8)),
	5817 => std_logic_vector(to_unsigned(42, 8)),
	5818 => std_logic_vector(to_unsigned(41, 8)),
	5819 => std_logic_vector(to_unsigned(42, 8)),
	5820 => std_logic_vector(to_unsigned(41, 8)),
	5821 => std_logic_vector(to_unsigned(42, 8)),
	5822 => std_logic_vector(to_unsigned(41, 8)),
	5823 => std_logic_vector(to_unsigned(42, 8)),
	5824 => std_logic_vector(to_unsigned(42, 8)),
	5825 => std_logic_vector(to_unsigned(42, 8)),
	5826 => std_logic_vector(to_unsigned(41, 8)),
	5827 => std_logic_vector(to_unsigned(42, 8)),
	5828 => std_logic_vector(to_unsigned(42, 8)),
	5829 => std_logic_vector(to_unsigned(41, 8)),
	5830 => std_logic_vector(to_unsigned(42, 8)),
	5831 => std_logic_vector(to_unsigned(41, 8)),
	5832 => std_logic_vector(to_unsigned(41, 8)),
	5833 => std_logic_vector(to_unsigned(41, 8)),
	5834 => std_logic_vector(to_unsigned(42, 8)),
	5835 => std_logic_vector(to_unsigned(42, 8)),
	5836 => std_logic_vector(to_unsigned(42, 8)),
	5837 => std_logic_vector(to_unsigned(41, 8)),
	5838 => std_logic_vector(to_unsigned(41, 8)),
	5839 => std_logic_vector(to_unsigned(42, 8)),
	5840 => std_logic_vector(to_unsigned(42, 8)),
	5841 => std_logic_vector(to_unsigned(41, 8)),
	5842 => std_logic_vector(to_unsigned(42, 8)),
	5843 => std_logic_vector(to_unsigned(42, 8)),
	5844 => std_logic_vector(to_unsigned(42, 8)),
	5845 => std_logic_vector(to_unsigned(42, 8)),
	5846 => std_logic_vector(to_unsigned(42, 8)),
	5847 => std_logic_vector(to_unsigned(41, 8)),
	5848 => std_logic_vector(to_unsigned(41, 8)),
	5849 => std_logic_vector(to_unsigned(41, 8)),
	5850 => std_logic_vector(to_unsigned(41, 8)),
	5851 => std_logic_vector(to_unsigned(42, 8)),
	5852 => std_logic_vector(to_unsigned(42, 8)),
	5853 => std_logic_vector(to_unsigned(42, 8)),
	5854 => std_logic_vector(to_unsigned(41, 8)),
	5855 => std_logic_vector(to_unsigned(41, 8)),
	5856 => std_logic_vector(to_unsigned(41, 8)),
	5857 => std_logic_vector(to_unsigned(42, 8)),
	5858 => std_logic_vector(to_unsigned(42, 8)),
	5859 => std_logic_vector(to_unsigned(42, 8)),
	5860 => std_logic_vector(to_unsigned(42, 8)),
	5861 => std_logic_vector(to_unsigned(41, 8)),
	5862 => std_logic_vector(to_unsigned(41, 8)),
	5863 => std_logic_vector(to_unsigned(42, 8)),
	5864 => std_logic_vector(to_unsigned(42, 8)),
	5865 => std_logic_vector(to_unsigned(41, 8)),
	5866 => std_logic_vector(to_unsigned(42, 8)),
	5867 => std_logic_vector(to_unsigned(42, 8)),
	5868 => std_logic_vector(to_unsigned(42, 8)),
	5869 => std_logic_vector(to_unsigned(42, 8)),
	5870 => std_logic_vector(to_unsigned(41, 8)),
	5871 => std_logic_vector(to_unsigned(42, 8)),
	5872 => std_logic_vector(to_unsigned(41, 8)),
	5873 => std_logic_vector(to_unsigned(42, 8)),
	5874 => std_logic_vector(to_unsigned(42, 8)),
	5875 => std_logic_vector(to_unsigned(42, 8)),
	5876 => std_logic_vector(to_unsigned(42, 8)),
	5877 => std_logic_vector(to_unsigned(41, 8)),
	5878 => std_logic_vector(to_unsigned(41, 8)),
	5879 => std_logic_vector(to_unsigned(42, 8)),
	5880 => std_logic_vector(to_unsigned(41, 8)),
	5881 => std_logic_vector(to_unsigned(41, 8)),
	5882 => std_logic_vector(to_unsigned(41, 8)),
	5883 => std_logic_vector(to_unsigned(41, 8)),
	5884 => std_logic_vector(to_unsigned(41, 8)),
	5885 => std_logic_vector(to_unsigned(42, 8)),
	5886 => std_logic_vector(to_unsigned(42, 8)),
	5887 => std_logic_vector(to_unsigned(42, 8)),
	5888 => std_logic_vector(to_unsigned(42, 8)),
	5889 => std_logic_vector(to_unsigned(41, 8)),
	5890 => std_logic_vector(to_unsigned(42, 8)),
	5891 => std_logic_vector(to_unsigned(42, 8)),
	5892 => std_logic_vector(to_unsigned(41, 8)),
	5893 => std_logic_vector(to_unsigned(41, 8)),
	5894 => std_logic_vector(to_unsigned(42, 8)),
	5895 => std_logic_vector(to_unsigned(42, 8)),
	5896 => std_logic_vector(to_unsigned(41, 8)),
	5897 => std_logic_vector(to_unsigned(41, 8)),
	5898 => std_logic_vector(to_unsigned(42, 8)),
	5899 => std_logic_vector(to_unsigned(41, 8)),
	5900 => std_logic_vector(to_unsigned(41, 8)),
	5901 => std_logic_vector(to_unsigned(41, 8)),
	5902 => std_logic_vector(to_unsigned(42, 8)),
	5903 => std_logic_vector(to_unsigned(42, 8)),
	5904 => std_logic_vector(to_unsigned(41, 8)),
	5905 => std_logic_vector(to_unsigned(41, 8)),
	5906 => std_logic_vector(to_unsigned(41, 8)),
	5907 => std_logic_vector(to_unsigned(41, 8)),
	5908 => std_logic_vector(to_unsigned(41, 8)),
	5909 => std_logic_vector(to_unsigned(41, 8)),
	5910 => std_logic_vector(to_unsigned(41, 8)),
	5911 => std_logic_vector(to_unsigned(42, 8)),
	5912 => std_logic_vector(to_unsigned(42, 8)),
	5913 => std_logic_vector(to_unsigned(41, 8)),
	5914 => std_logic_vector(to_unsigned(42, 8)),
	5915 => std_logic_vector(to_unsigned(42, 8)),
	5916 => std_logic_vector(to_unsigned(41, 8)),
	5917 => std_logic_vector(to_unsigned(42, 8)),
	5918 => std_logic_vector(to_unsigned(41, 8)),
	5919 => std_logic_vector(to_unsigned(41, 8)),
	5920 => std_logic_vector(to_unsigned(41, 8)),
	5921 => std_logic_vector(to_unsigned(41, 8)),
	5922 => std_logic_vector(to_unsigned(41, 8)),
	5923 => std_logic_vector(to_unsigned(41, 8)),
	5924 => std_logic_vector(to_unsigned(41, 8)),
	5925 => std_logic_vector(to_unsigned(41, 8)),
	5926 => std_logic_vector(to_unsigned(42, 8)),
	5927 => std_logic_vector(to_unsigned(42, 8)),
	5928 => std_logic_vector(to_unsigned(41, 8)),
	5929 => std_logic_vector(to_unsigned(41, 8)),
	5930 => std_logic_vector(to_unsigned(42, 8)),
	5931 => std_logic_vector(to_unsigned(41, 8)),
	5932 => std_logic_vector(to_unsigned(41, 8)),
	5933 => std_logic_vector(to_unsigned(41, 8)),
	5934 => std_logic_vector(to_unsigned(41, 8)),
	5935 => std_logic_vector(to_unsigned(42, 8)),
	5936 => std_logic_vector(to_unsigned(41, 8)),
	5937 => std_logic_vector(to_unsigned(42, 8)),
	5938 => std_logic_vector(to_unsigned(41, 8)),
	5939 => std_logic_vector(to_unsigned(42, 8)),
	5940 => std_logic_vector(to_unsigned(41, 8)),
	5941 => std_logic_vector(to_unsigned(41, 8)),
	5942 => std_logic_vector(to_unsigned(41, 8)),
	5943 => std_logic_vector(to_unsigned(42, 8)),
	5944 => std_logic_vector(to_unsigned(41, 8)),
	5945 => std_logic_vector(to_unsigned(42, 8)),
	5946 => std_logic_vector(to_unsigned(41, 8)),
	5947 => std_logic_vector(to_unsigned(41, 8)),
	5948 => std_logic_vector(to_unsigned(41, 8)),
	5949 => std_logic_vector(to_unsigned(42, 8)),
	5950 => std_logic_vector(to_unsigned(42, 8)),
	5951 => std_logic_vector(to_unsigned(42, 8)),
	5952 => std_logic_vector(to_unsigned(42, 8)),
	5953 => std_logic_vector(to_unsigned(41, 8)),
	5954 => std_logic_vector(to_unsigned(42, 8)),
	5955 => std_logic_vector(to_unsigned(42, 8)),
	5956 => std_logic_vector(to_unsigned(42, 8)),
	5957 => std_logic_vector(to_unsigned(42, 8)),
	5958 => std_logic_vector(to_unsigned(42, 8)),
	5959 => std_logic_vector(to_unsigned(42, 8)),
	5960 => std_logic_vector(to_unsigned(42, 8)),
	5961 => std_logic_vector(to_unsigned(41, 8)),
	5962 => std_logic_vector(to_unsigned(41, 8)),
	5963 => std_logic_vector(to_unsigned(41, 8)),
	5964 => std_logic_vector(to_unsigned(42, 8)),
	5965 => std_logic_vector(to_unsigned(41, 8)),
	5966 => std_logic_vector(to_unsigned(41, 8)),
	5967 => std_logic_vector(to_unsigned(42, 8)),
	5968 => std_logic_vector(to_unsigned(42, 8)),
	5969 => std_logic_vector(to_unsigned(42, 8)),
	5970 => std_logic_vector(to_unsigned(41, 8)),
	5971 => std_logic_vector(to_unsigned(41, 8)),
	5972 => std_logic_vector(to_unsigned(42, 8)),
	5973 => std_logic_vector(to_unsigned(42, 8)),
	5974 => std_logic_vector(to_unsigned(42, 8)),
	5975 => std_logic_vector(to_unsigned(41, 8)),
	5976 => std_logic_vector(to_unsigned(42, 8)),
	5977 => std_logic_vector(to_unsigned(41, 8)),
	5978 => std_logic_vector(to_unsigned(42, 8)),
	5979 => std_logic_vector(to_unsigned(42, 8)),
	5980 => std_logic_vector(to_unsigned(42, 8)),
	5981 => std_logic_vector(to_unsigned(41, 8)),
	5982 => std_logic_vector(to_unsigned(41, 8)),
	5983 => std_logic_vector(to_unsigned(42, 8)),
	5984 => std_logic_vector(to_unsigned(41, 8)),
	5985 => std_logic_vector(to_unsigned(42, 8)),
	5986 => std_logic_vector(to_unsigned(41, 8)),
	5987 => std_logic_vector(to_unsigned(42, 8)),
	5988 => std_logic_vector(to_unsigned(41, 8)),
	5989 => std_logic_vector(to_unsigned(42, 8)),
	5990 => std_logic_vector(to_unsigned(42, 8)),
	5991 => std_logic_vector(to_unsigned(41, 8)),
	5992 => std_logic_vector(to_unsigned(42, 8)),
	5993 => std_logic_vector(to_unsigned(42, 8)),
	5994 => std_logic_vector(to_unsigned(41, 8)),
	5995 => std_logic_vector(to_unsigned(41, 8)),
	5996 => std_logic_vector(to_unsigned(41, 8)),
	5997 => std_logic_vector(to_unsigned(41, 8)),
	5998 => std_logic_vector(to_unsigned(41, 8)),
	5999 => std_logic_vector(to_unsigned(41, 8)),
	6000 => std_logic_vector(to_unsigned(41, 8)),
	6001 => std_logic_vector(to_unsigned(42, 8)),
	6002 => std_logic_vector(to_unsigned(42, 8)),
	6003 => std_logic_vector(to_unsigned(41, 8)),
	6004 => std_logic_vector(to_unsigned(41, 8)),
	6005 => std_logic_vector(to_unsigned(42, 8)),
	6006 => std_logic_vector(to_unsigned(41, 8)),
	6007 => std_logic_vector(to_unsigned(42, 8)),
	6008 => std_logic_vector(to_unsigned(42, 8)),
	6009 => std_logic_vector(to_unsigned(42, 8)),
	6010 => std_logic_vector(to_unsigned(42, 8)),
	6011 => std_logic_vector(to_unsigned(42, 8)),
	6012 => std_logic_vector(to_unsigned(41, 8)),
	6013 => std_logic_vector(to_unsigned(41, 8)),
	6014 => std_logic_vector(to_unsigned(42, 8)),
	6015 => std_logic_vector(to_unsigned(42, 8)),
	6016 => std_logic_vector(to_unsigned(41, 8)),
	6017 => std_logic_vector(to_unsigned(41, 8)),
	6018 => std_logic_vector(to_unsigned(41, 8)),
	6019 => std_logic_vector(to_unsigned(42, 8)),
	6020 => std_logic_vector(to_unsigned(42, 8)),
	6021 => std_logic_vector(to_unsigned(41, 8)),
	6022 => std_logic_vector(to_unsigned(42, 8)),
	6023 => std_logic_vector(to_unsigned(41, 8)),
	6024 => std_logic_vector(to_unsigned(41, 8)),
	6025 => std_logic_vector(to_unsigned(42, 8)),
	6026 => std_logic_vector(to_unsigned(41, 8)),
	6027 => std_logic_vector(to_unsigned(42, 8)),
	6028 => std_logic_vector(to_unsigned(41, 8)),
	6029 => std_logic_vector(to_unsigned(42, 8)),
	6030 => std_logic_vector(to_unsigned(42, 8)),
	6031 => std_logic_vector(to_unsigned(42, 8)),
	6032 => std_logic_vector(to_unsigned(41, 8)),
	6033 => std_logic_vector(to_unsigned(41, 8)),
	6034 => std_logic_vector(to_unsigned(41, 8)),
	6035 => std_logic_vector(to_unsigned(41, 8)),
	6036 => std_logic_vector(to_unsigned(42, 8)),
	6037 => std_logic_vector(to_unsigned(41, 8)),
	6038 => std_logic_vector(to_unsigned(41, 8)),
	6039 => std_logic_vector(to_unsigned(42, 8)),
	6040 => std_logic_vector(to_unsigned(42, 8)),
	6041 => std_logic_vector(to_unsigned(41, 8)),
	6042 => std_logic_vector(to_unsigned(41, 8)),
	6043 => std_logic_vector(to_unsigned(42, 8)),
	6044 => std_logic_vector(to_unsigned(41, 8)),
	6045 => std_logic_vector(to_unsigned(41, 8)),
	6046 => std_logic_vector(to_unsigned(42, 8)),
	6047 => std_logic_vector(to_unsigned(41, 8)),
	6048 => std_logic_vector(to_unsigned(41, 8)),
	6049 => std_logic_vector(to_unsigned(41, 8)),
	6050 => std_logic_vector(to_unsigned(42, 8)),
	6051 => std_logic_vector(to_unsigned(42, 8)),
	6052 => std_logic_vector(to_unsigned(41, 8)),
	6053 => std_logic_vector(to_unsigned(42, 8)),
	6054 => std_logic_vector(to_unsigned(42, 8)),
	6055 => std_logic_vector(to_unsigned(41, 8)),
	6056 => std_logic_vector(to_unsigned(41, 8)),
	6057 => std_logic_vector(to_unsigned(42, 8)),
	6058 => std_logic_vector(to_unsigned(41, 8)),
	6059 => std_logic_vector(to_unsigned(41, 8)),
	6060 => std_logic_vector(to_unsigned(41, 8)),
	6061 => std_logic_vector(to_unsigned(42, 8)),
	6062 => std_logic_vector(to_unsigned(42, 8)),
	6063 => std_logic_vector(to_unsigned(41, 8)),
	6064 => std_logic_vector(to_unsigned(42, 8)),
	6065 => std_logic_vector(to_unsigned(41, 8)),
	6066 => std_logic_vector(to_unsigned(41, 8)),
	6067 => std_logic_vector(to_unsigned(42, 8)),
	6068 => std_logic_vector(to_unsigned(41, 8)),
	6069 => std_logic_vector(to_unsigned(41, 8)),
	6070 => std_logic_vector(to_unsigned(41, 8)),
	6071 => std_logic_vector(to_unsigned(42, 8)),
	6072 => std_logic_vector(to_unsigned(41, 8)),
	6073 => std_logic_vector(to_unsigned(42, 8)),
	6074 => std_logic_vector(to_unsigned(42, 8)),
	6075 => std_logic_vector(to_unsigned(42, 8)),
	6076 => std_logic_vector(to_unsigned(42, 8)),
	6077 => std_logic_vector(to_unsigned(41, 8)),
	6078 => std_logic_vector(to_unsigned(41, 8)),
	6079 => std_logic_vector(to_unsigned(41, 8)),
	6080 => std_logic_vector(to_unsigned(42, 8)),
	6081 => std_logic_vector(to_unsigned(42, 8)),
	6082 => std_logic_vector(to_unsigned(41, 8)),
	6083 => std_logic_vector(to_unsigned(41, 8)),
	6084 => std_logic_vector(to_unsigned(42, 8)),
	6085 => std_logic_vector(to_unsigned(42, 8)),
	6086 => std_logic_vector(to_unsigned(42, 8)),
	6087 => std_logic_vector(to_unsigned(41, 8)),
	6088 => std_logic_vector(to_unsigned(42, 8)),
	6089 => std_logic_vector(to_unsigned(42, 8)),
	6090 => std_logic_vector(to_unsigned(42, 8)),
	6091 => std_logic_vector(to_unsigned(41, 8)),
	6092 => std_logic_vector(to_unsigned(42, 8)),
	6093 => std_logic_vector(to_unsigned(41, 8)),
	6094 => std_logic_vector(to_unsigned(41, 8)),
	6095 => std_logic_vector(to_unsigned(41, 8)),
	6096 => std_logic_vector(to_unsigned(41, 8)),
	6097 => std_logic_vector(to_unsigned(41, 8)),
	6098 => std_logic_vector(to_unsigned(42, 8)),
	6099 => std_logic_vector(to_unsigned(41, 8)),
	6100 => std_logic_vector(to_unsigned(42, 8)),
	6101 => std_logic_vector(to_unsigned(41, 8)),
	6102 => std_logic_vector(to_unsigned(41, 8)),
	6103 => std_logic_vector(to_unsigned(41, 8)),
	6104 => std_logic_vector(to_unsigned(41, 8)),
	6105 => std_logic_vector(to_unsigned(42, 8)),
	6106 => std_logic_vector(to_unsigned(41, 8)),
	6107 => std_logic_vector(to_unsigned(41, 8)),
	6108 => std_logic_vector(to_unsigned(41, 8)),
	6109 => std_logic_vector(to_unsigned(41, 8)),
	6110 => std_logic_vector(to_unsigned(41, 8)),
	6111 => std_logic_vector(to_unsigned(41, 8)),
	6112 => std_logic_vector(to_unsigned(42, 8)),
	6113 => std_logic_vector(to_unsigned(42, 8)),
	6114 => std_logic_vector(to_unsigned(42, 8)),
	6115 => std_logic_vector(to_unsigned(41, 8)),
	6116 => std_logic_vector(to_unsigned(42, 8)),
	6117 => std_logic_vector(to_unsigned(41, 8)),
	6118 => std_logic_vector(to_unsigned(42, 8)),
	6119 => std_logic_vector(to_unsigned(41, 8)),
	6120 => std_logic_vector(to_unsigned(41, 8)),
	6121 => std_logic_vector(to_unsigned(42, 8)),
	6122 => std_logic_vector(to_unsigned(41, 8)),
	6123 => std_logic_vector(to_unsigned(41, 8)),
	6124 => std_logic_vector(to_unsigned(41, 8)),
	6125 => std_logic_vector(to_unsigned(42, 8)),
	6126 => std_logic_vector(to_unsigned(41, 8)),
	6127 => std_logic_vector(to_unsigned(42, 8)),
	6128 => std_logic_vector(to_unsigned(42, 8)),
	6129 => std_logic_vector(to_unsigned(42, 8)),
	6130 => std_logic_vector(to_unsigned(41, 8)),
	6131 => std_logic_vector(to_unsigned(42, 8)),
	6132 => std_logic_vector(to_unsigned(41, 8)),
	6133 => std_logic_vector(to_unsigned(42, 8)),
	6134 => std_logic_vector(to_unsigned(42, 8)),
	6135 => std_logic_vector(to_unsigned(42, 8)),
	6136 => std_logic_vector(to_unsigned(42, 8)),
	6137 => std_logic_vector(to_unsigned(41, 8)),
	6138 => std_logic_vector(to_unsigned(41, 8)),
	6139 => std_logic_vector(to_unsigned(41, 8)),
	6140 => std_logic_vector(to_unsigned(41, 8)),
	6141 => std_logic_vector(to_unsigned(42, 8)),
	6142 => std_logic_vector(to_unsigned(42, 8)),
	6143 => std_logic_vector(to_unsigned(41, 8)),
	6144 => std_logic_vector(to_unsigned(42, 8)),
	6145 => std_logic_vector(to_unsigned(41, 8)),
	6146 => std_logic_vector(to_unsigned(41, 8)),
	6147 => std_logic_vector(to_unsigned(41, 8)),
	6148 => std_logic_vector(to_unsigned(41, 8)),
	6149 => std_logic_vector(to_unsigned(41, 8)),
	6150 => std_logic_vector(to_unsigned(41, 8)),
	6151 => std_logic_vector(to_unsigned(42, 8)),
	6152 => std_logic_vector(to_unsigned(41, 8)),
	6153 => std_logic_vector(to_unsigned(42, 8)),
	6154 => std_logic_vector(to_unsigned(42, 8)),
	6155 => std_logic_vector(to_unsigned(42, 8)),
	6156 => std_logic_vector(to_unsigned(41, 8)),
	6157 => std_logic_vector(to_unsigned(41, 8)),
	6158 => std_logic_vector(to_unsigned(42, 8)),
	6159 => std_logic_vector(to_unsigned(41, 8)),
	6160 => std_logic_vector(to_unsigned(42, 8)),
	6161 => std_logic_vector(to_unsigned(41, 8)),
	6162 => std_logic_vector(to_unsigned(41, 8)),
	6163 => std_logic_vector(to_unsigned(42, 8)),
	6164 => std_logic_vector(to_unsigned(41, 8)),
	6165 => std_logic_vector(to_unsigned(42, 8)),
	6166 => std_logic_vector(to_unsigned(41, 8)),
	6167 => std_logic_vector(to_unsigned(42, 8)),
	6168 => std_logic_vector(to_unsigned(41, 8)),
	6169 => std_logic_vector(to_unsigned(42, 8)),
	6170 => std_logic_vector(to_unsigned(41, 8)),
	6171 => std_logic_vector(to_unsigned(42, 8)),
	6172 => std_logic_vector(to_unsigned(42, 8)),
	6173 => std_logic_vector(to_unsigned(41, 8)),
	6174 => std_logic_vector(to_unsigned(41, 8)),
	6175 => std_logic_vector(to_unsigned(41, 8)),
	6176 => std_logic_vector(to_unsigned(42, 8)),
	6177 => std_logic_vector(to_unsigned(41, 8)),
	6178 => std_logic_vector(to_unsigned(41, 8)),
	6179 => std_logic_vector(to_unsigned(42, 8)),
	6180 => std_logic_vector(to_unsigned(42, 8)),
	6181 => std_logic_vector(to_unsigned(41, 8)),
	6182 => std_logic_vector(to_unsigned(42, 8)),
	6183 => std_logic_vector(to_unsigned(41, 8)),
	6184 => std_logic_vector(to_unsigned(42, 8)),
	6185 => std_logic_vector(to_unsigned(42, 8)),
	6186 => std_logic_vector(to_unsigned(41, 8)),
	6187 => std_logic_vector(to_unsigned(42, 8)),
	6188 => std_logic_vector(to_unsigned(42, 8)),
	6189 => std_logic_vector(to_unsigned(42, 8)),
	6190 => std_logic_vector(to_unsigned(42, 8)),
	6191 => std_logic_vector(to_unsigned(41, 8)),
	6192 => std_logic_vector(to_unsigned(42, 8)),
	6193 => std_logic_vector(to_unsigned(41, 8)),
	6194 => std_logic_vector(to_unsigned(42, 8)),
	6195 => std_logic_vector(to_unsigned(41, 8)),
	6196 => std_logic_vector(to_unsigned(41, 8)),
	6197 => std_logic_vector(to_unsigned(42, 8)),
	6198 => std_logic_vector(to_unsigned(42, 8)),
	6199 => std_logic_vector(to_unsigned(42, 8)),
	6200 => std_logic_vector(to_unsigned(42, 8)),
	6201 => std_logic_vector(to_unsigned(42, 8)),
	6202 => std_logic_vector(to_unsigned(42, 8)),
	6203 => std_logic_vector(to_unsigned(42, 8)),
	6204 => std_logic_vector(to_unsigned(41, 8)),
	6205 => std_logic_vector(to_unsigned(41, 8)),
	6206 => std_logic_vector(to_unsigned(42, 8)),
	6207 => std_logic_vector(to_unsigned(42, 8)),
	6208 => std_logic_vector(to_unsigned(41, 8)),
	6209 => std_logic_vector(to_unsigned(41, 8)),
	6210 => std_logic_vector(to_unsigned(42, 8)),
	6211 => std_logic_vector(to_unsigned(42, 8)),
	6212 => std_logic_vector(to_unsigned(42, 8)),
	6213 => std_logic_vector(to_unsigned(41, 8)),
	6214 => std_logic_vector(to_unsigned(42, 8)),
	6215 => std_logic_vector(to_unsigned(41, 8)),
	6216 => std_logic_vector(to_unsigned(41, 8)),
	6217 => std_logic_vector(to_unsigned(41, 8)),
	6218 => std_logic_vector(to_unsigned(41, 8)),
	6219 => std_logic_vector(to_unsigned(42, 8)),
	6220 => std_logic_vector(to_unsigned(41, 8)),
	6221 => std_logic_vector(to_unsigned(42, 8)),
	6222 => std_logic_vector(to_unsigned(41, 8)),
	6223 => std_logic_vector(to_unsigned(41, 8)),
	6224 => std_logic_vector(to_unsigned(41, 8)),
	6225 => std_logic_vector(to_unsigned(42, 8)),
	6226 => std_logic_vector(to_unsigned(41, 8)),
	6227 => std_logic_vector(to_unsigned(42, 8)),
	6228 => std_logic_vector(to_unsigned(42, 8)),
	6229 => std_logic_vector(to_unsigned(41, 8)),
	6230 => std_logic_vector(to_unsigned(41, 8)),
	6231 => std_logic_vector(to_unsigned(42, 8)),
	6232 => std_logic_vector(to_unsigned(42, 8)),
	6233 => std_logic_vector(to_unsigned(41, 8)),
	6234 => std_logic_vector(to_unsigned(42, 8)),
	6235 => std_logic_vector(to_unsigned(41, 8)),
	6236 => std_logic_vector(to_unsigned(41, 8)),
	6237 => std_logic_vector(to_unsigned(42, 8)),
	6238 => std_logic_vector(to_unsigned(41, 8)),
	6239 => std_logic_vector(to_unsigned(42, 8)),
	6240 => std_logic_vector(to_unsigned(42, 8)),
	6241 => std_logic_vector(to_unsigned(42, 8)),
	6242 => std_logic_vector(to_unsigned(42, 8)),
	6243 => std_logic_vector(to_unsigned(41, 8)),
	6244 => std_logic_vector(to_unsigned(41, 8)),
	6245 => std_logic_vector(to_unsigned(42, 8)),
	6246 => std_logic_vector(to_unsigned(42, 8)),
	6247 => std_logic_vector(to_unsigned(41, 8)),
	6248 => std_logic_vector(to_unsigned(41, 8)),
	6249 => std_logic_vector(to_unsigned(42, 8)),
	6250 => std_logic_vector(to_unsigned(42, 8)),
	6251 => std_logic_vector(to_unsigned(41, 8)),
	6252 => std_logic_vector(to_unsigned(42, 8)),
	6253 => std_logic_vector(to_unsigned(42, 8)),
	6254 => std_logic_vector(to_unsigned(41, 8)),
	6255 => std_logic_vector(to_unsigned(42, 8)),
	6256 => std_logic_vector(to_unsigned(42, 8)),
	6257 => std_logic_vector(to_unsigned(42, 8)),
	6258 => std_logic_vector(to_unsigned(42, 8)),
	6259 => std_logic_vector(to_unsigned(42, 8)),
	6260 => std_logic_vector(to_unsigned(41, 8)),
	6261 => std_logic_vector(to_unsigned(42, 8)),
	6262 => std_logic_vector(to_unsigned(41, 8)),
	6263 => std_logic_vector(to_unsigned(42, 8)),
	6264 => std_logic_vector(to_unsigned(42, 8)),
	6265 => std_logic_vector(to_unsigned(42, 8)),
	6266 => std_logic_vector(to_unsigned(41, 8)),
	6267 => std_logic_vector(to_unsigned(42, 8)),
	6268 => std_logic_vector(to_unsigned(42, 8)),
	6269 => std_logic_vector(to_unsigned(42, 8)),
	6270 => std_logic_vector(to_unsigned(42, 8)),
	6271 => std_logic_vector(to_unsigned(42, 8)),
	6272 => std_logic_vector(to_unsigned(41, 8)),
	6273 => std_logic_vector(to_unsigned(42, 8)),
	6274 => std_logic_vector(to_unsigned(41, 8)),
	6275 => std_logic_vector(to_unsigned(42, 8)),
	6276 => std_logic_vector(to_unsigned(42, 8)),
	6277 => std_logic_vector(to_unsigned(42, 8)),
	6278 => std_logic_vector(to_unsigned(41, 8)),
	6279 => std_logic_vector(to_unsigned(42, 8)),
	6280 => std_logic_vector(to_unsigned(41, 8)),
	6281 => std_logic_vector(to_unsigned(42, 8)),
	6282 => std_logic_vector(to_unsigned(42, 8)),
	6283 => std_logic_vector(to_unsigned(42, 8)),
	6284 => std_logic_vector(to_unsigned(41, 8)),
	6285 => std_logic_vector(to_unsigned(42, 8)),
	6286 => std_logic_vector(to_unsigned(41, 8)),
	6287 => std_logic_vector(to_unsigned(42, 8)),
	6288 => std_logic_vector(to_unsigned(42, 8)),
	6289 => std_logic_vector(to_unsigned(42, 8)),
	6290 => std_logic_vector(to_unsigned(41, 8)),
	6291 => std_logic_vector(to_unsigned(41, 8)),
	6292 => std_logic_vector(to_unsigned(42, 8)),
	6293 => std_logic_vector(to_unsigned(41, 8)),
	6294 => std_logic_vector(to_unsigned(41, 8)),
	6295 => std_logic_vector(to_unsigned(42, 8)),
	6296 => std_logic_vector(to_unsigned(42, 8)),
	6297 => std_logic_vector(to_unsigned(41, 8)),
	6298 => std_logic_vector(to_unsigned(41, 8)),
	6299 => std_logic_vector(to_unsigned(42, 8)),
	6300 => std_logic_vector(to_unsigned(42, 8)),
	6301 => std_logic_vector(to_unsigned(41, 8)),
	6302 => std_logic_vector(to_unsigned(42, 8)),
	6303 => std_logic_vector(to_unsigned(42, 8)),
	6304 => std_logic_vector(to_unsigned(41, 8)),
	6305 => std_logic_vector(to_unsigned(42, 8)),
	6306 => std_logic_vector(to_unsigned(42, 8)),
	6307 => std_logic_vector(to_unsigned(42, 8)),
	6308 => std_logic_vector(to_unsigned(42, 8)),
	6309 => std_logic_vector(to_unsigned(42, 8)),
	6310 => std_logic_vector(to_unsigned(41, 8)),
	6311 => std_logic_vector(to_unsigned(42, 8)),
	6312 => std_logic_vector(to_unsigned(41, 8)),
	6313 => std_logic_vector(to_unsigned(42, 8)),
	6314 => std_logic_vector(to_unsigned(41, 8)),
	6315 => std_logic_vector(to_unsigned(41, 8)),
	6316 => std_logic_vector(to_unsigned(42, 8)),
	6317 => std_logic_vector(to_unsigned(42, 8)),
	6318 => std_logic_vector(to_unsigned(42, 8)),
	6319 => std_logic_vector(to_unsigned(41, 8)),
	6320 => std_logic_vector(to_unsigned(42, 8)),
	6321 => std_logic_vector(to_unsigned(42, 8)),
	6322 => std_logic_vector(to_unsigned(41, 8)),
	6323 => std_logic_vector(to_unsigned(41, 8)),
	6324 => std_logic_vector(to_unsigned(42, 8)),
	6325 => std_logic_vector(to_unsigned(41, 8)),
	6326 => std_logic_vector(to_unsigned(42, 8)),
	6327 => std_logic_vector(to_unsigned(42, 8)),
	6328 => std_logic_vector(to_unsigned(42, 8)),
	6329 => std_logic_vector(to_unsigned(42, 8)),
	6330 => std_logic_vector(to_unsigned(41, 8)),
	6331 => std_logic_vector(to_unsigned(41, 8)),
	6332 => std_logic_vector(to_unsigned(42, 8)),
	6333 => std_logic_vector(to_unsigned(41, 8)),
	6334 => std_logic_vector(to_unsigned(42, 8)),
	6335 => std_logic_vector(to_unsigned(42, 8)),
	6336 => std_logic_vector(to_unsigned(42, 8)),
	6337 => std_logic_vector(to_unsigned(41, 8)),
	6338 => std_logic_vector(to_unsigned(41, 8)),
	6339 => std_logic_vector(to_unsigned(41, 8)),
	6340 => std_logic_vector(to_unsigned(41, 8)),
	6341 => std_logic_vector(to_unsigned(41, 8)),
	6342 => std_logic_vector(to_unsigned(42, 8)),
	6343 => std_logic_vector(to_unsigned(42, 8)),
	6344 => std_logic_vector(to_unsigned(42, 8)),
	6345 => std_logic_vector(to_unsigned(42, 8)),
	6346 => std_logic_vector(to_unsigned(42, 8)),
	6347 => std_logic_vector(to_unsigned(42, 8)),
	6348 => std_logic_vector(to_unsigned(42, 8)),
	6349 => std_logic_vector(to_unsigned(41, 8)),
	6350 => std_logic_vector(to_unsigned(41, 8)),
	6351 => std_logic_vector(to_unsigned(41, 8)),
	6352 => std_logic_vector(to_unsigned(41, 8)),
	6353 => std_logic_vector(to_unsigned(42, 8)),
	6354 => std_logic_vector(to_unsigned(42, 8)),
	6355 => std_logic_vector(to_unsigned(41, 8)),
	6356 => std_logic_vector(to_unsigned(41, 8)),
	6357 => std_logic_vector(to_unsigned(41, 8)),
	6358 => std_logic_vector(to_unsigned(41, 8)),
	6359 => std_logic_vector(to_unsigned(41, 8)),
	6360 => std_logic_vector(to_unsigned(42, 8)),
	6361 => std_logic_vector(to_unsigned(41, 8)),
	6362 => std_logic_vector(to_unsigned(41, 8)),
	6363 => std_logic_vector(to_unsigned(42, 8)),
	6364 => std_logic_vector(to_unsigned(41, 8)),
	6365 => std_logic_vector(to_unsigned(41, 8)),
	6366 => std_logic_vector(to_unsigned(41, 8)),
	6367 => std_logic_vector(to_unsigned(42, 8)),
	6368 => std_logic_vector(to_unsigned(41, 8)),
	6369 => std_logic_vector(to_unsigned(41, 8)),
	6370 => std_logic_vector(to_unsigned(42, 8)),
	6371 => std_logic_vector(to_unsigned(41, 8)),
	6372 => std_logic_vector(to_unsigned(41, 8)),
	6373 => std_logic_vector(to_unsigned(41, 8)),
	6374 => std_logic_vector(to_unsigned(41, 8)),
	6375 => std_logic_vector(to_unsigned(41, 8)),
	6376 => std_logic_vector(to_unsigned(41, 8)),
	6377 => std_logic_vector(to_unsigned(42, 8)),
	6378 => std_logic_vector(to_unsigned(42, 8)),
	6379 => std_logic_vector(to_unsigned(41, 8)),
	6380 => std_logic_vector(to_unsigned(42, 8)),
	6381 => std_logic_vector(to_unsigned(42, 8)),
	6382 => std_logic_vector(to_unsigned(42, 8)),
	6383 => std_logic_vector(to_unsigned(42, 8)),
	6384 => std_logic_vector(to_unsigned(41, 8)),
	6385 => std_logic_vector(to_unsigned(41, 8)),
	6386 => std_logic_vector(to_unsigned(41, 8)),
	6387 => std_logic_vector(to_unsigned(42, 8)),
	6388 => std_logic_vector(to_unsigned(41, 8)),
	6389 => std_logic_vector(to_unsigned(42, 8)),
	6390 => std_logic_vector(to_unsigned(41, 8)),
	6391 => std_logic_vector(to_unsigned(41, 8)),
	6392 => std_logic_vector(to_unsigned(41, 8)),
	6393 => std_logic_vector(to_unsigned(42, 8)),
	6394 => std_logic_vector(to_unsigned(42, 8)),
	6395 => std_logic_vector(to_unsigned(42, 8)),
	6396 => std_logic_vector(to_unsigned(42, 8)),
	6397 => std_logic_vector(to_unsigned(42, 8)),
	6398 => std_logic_vector(to_unsigned(42, 8)),
	6399 => std_logic_vector(to_unsigned(41, 8)),
	6400 => std_logic_vector(to_unsigned(42, 8)),
	6401 => std_logic_vector(to_unsigned(41, 8)),
	6402 => std_logic_vector(to_unsigned(41, 8)),
	6403 => std_logic_vector(to_unsigned(41, 8)),
	6404 => std_logic_vector(to_unsigned(42, 8)),
	6405 => std_logic_vector(to_unsigned(42, 8)),
	6406 => std_logic_vector(to_unsigned(41, 8)),
	6407 => std_logic_vector(to_unsigned(42, 8)),
	6408 => std_logic_vector(to_unsigned(41, 8)),
	6409 => std_logic_vector(to_unsigned(42, 8)),
	6410 => std_logic_vector(to_unsigned(42, 8)),
	6411 => std_logic_vector(to_unsigned(42, 8)),
	6412 => std_logic_vector(to_unsigned(41, 8)),
	6413 => std_logic_vector(to_unsigned(42, 8)),
	6414 => std_logic_vector(to_unsigned(42, 8)),
	6415 => std_logic_vector(to_unsigned(42, 8)),
	6416 => std_logic_vector(to_unsigned(42, 8)),
	6417 => std_logic_vector(to_unsigned(42, 8)),
	6418 => std_logic_vector(to_unsigned(41, 8)),
	6419 => std_logic_vector(to_unsigned(41, 8)),
	6420 => std_logic_vector(to_unsigned(42, 8)),
	6421 => std_logic_vector(to_unsigned(41, 8)),
	6422 => std_logic_vector(to_unsigned(42, 8)),
	6423 => std_logic_vector(to_unsigned(42, 8)),
	6424 => std_logic_vector(to_unsigned(41, 8)),
	6425 => std_logic_vector(to_unsigned(42, 8)),
	6426 => std_logic_vector(to_unsigned(42, 8)),
	6427 => std_logic_vector(to_unsigned(41, 8)),
	6428 => std_logic_vector(to_unsigned(42, 8)),
	6429 => std_logic_vector(to_unsigned(42, 8)),
	6430 => std_logic_vector(to_unsigned(42, 8)),
	6431 => std_logic_vector(to_unsigned(41, 8)),
	6432 => std_logic_vector(to_unsigned(41, 8)),
	6433 => std_logic_vector(to_unsigned(41, 8)),
	6434 => std_logic_vector(to_unsigned(42, 8)),
	6435 => std_logic_vector(to_unsigned(42, 8)),
	6436 => std_logic_vector(to_unsigned(41, 8)),
	6437 => std_logic_vector(to_unsigned(42, 8)),
	6438 => std_logic_vector(to_unsigned(42, 8)),
	6439 => std_logic_vector(to_unsigned(42, 8)),
	6440 => std_logic_vector(to_unsigned(42, 8)),
	6441 => std_logic_vector(to_unsigned(42, 8)),
	6442 => std_logic_vector(to_unsigned(42, 8)),
	6443 => std_logic_vector(to_unsigned(41, 8)),
	6444 => std_logic_vector(to_unsigned(42, 8)),
	6445 => std_logic_vector(to_unsigned(41, 8)),
	6446 => std_logic_vector(to_unsigned(41, 8)),
	6447 => std_logic_vector(to_unsigned(42, 8)),
	6448 => std_logic_vector(to_unsigned(42, 8)),
	6449 => std_logic_vector(to_unsigned(41, 8)),
	6450 => std_logic_vector(to_unsigned(41, 8)),
	6451 => std_logic_vector(to_unsigned(42, 8)),
	6452 => std_logic_vector(to_unsigned(41, 8)),
	6453 => std_logic_vector(to_unsigned(41, 8)),
	6454 => std_logic_vector(to_unsigned(42, 8)),
	6455 => std_logic_vector(to_unsigned(41, 8)),
	6456 => std_logic_vector(to_unsigned(42, 8)),
	6457 => std_logic_vector(to_unsigned(41, 8)),
	6458 => std_logic_vector(to_unsigned(41, 8)),
	6459 => std_logic_vector(to_unsigned(42, 8)),
	6460 => std_logic_vector(to_unsigned(41, 8)),
	6461 => std_logic_vector(to_unsigned(42, 8)),
	6462 => std_logic_vector(to_unsigned(42, 8)),
	6463 => std_logic_vector(to_unsigned(42, 8)),
	6464 => std_logic_vector(to_unsigned(41, 8)),
	6465 => std_logic_vector(to_unsigned(42, 8)),
	6466 => std_logic_vector(to_unsigned(41, 8)),
	6467 => std_logic_vector(to_unsigned(41, 8)),
	6468 => std_logic_vector(to_unsigned(42, 8)),
	6469 => std_logic_vector(to_unsigned(41, 8)),
	6470 => std_logic_vector(to_unsigned(42, 8)),
	6471 => std_logic_vector(to_unsigned(42, 8)),
	6472 => std_logic_vector(to_unsigned(42, 8)),
	6473 => std_logic_vector(to_unsigned(42, 8)),
	6474 => std_logic_vector(to_unsigned(42, 8)),
	6475 => std_logic_vector(to_unsigned(42, 8)),
	6476 => std_logic_vector(to_unsigned(41, 8)),
	6477 => std_logic_vector(to_unsigned(41, 8)),
	6478 => std_logic_vector(to_unsigned(42, 8)),
	6479 => std_logic_vector(to_unsigned(41, 8)),
	6480 => std_logic_vector(to_unsigned(42, 8)),
	6481 => std_logic_vector(to_unsigned(42, 8)),
	6482 => std_logic_vector(to_unsigned(42, 8)),
	6483 => std_logic_vector(to_unsigned(42, 8)),
	6484 => std_logic_vector(to_unsigned(41, 8)),
	6485 => std_logic_vector(to_unsigned(42, 8)),
	6486 => std_logic_vector(to_unsigned(42, 8)),
	6487 => std_logic_vector(to_unsigned(42, 8)),
	6488 => std_logic_vector(to_unsigned(42, 8)),
	6489 => std_logic_vector(to_unsigned(42, 8)),
	6490 => std_logic_vector(to_unsigned(42, 8)),
	6491 => std_logic_vector(to_unsigned(42, 8)),
	6492 => std_logic_vector(to_unsigned(41, 8)),
	6493 => std_logic_vector(to_unsigned(41, 8)),
	6494 => std_logic_vector(to_unsigned(42, 8)),
	6495 => std_logic_vector(to_unsigned(41, 8)),
	6496 => std_logic_vector(to_unsigned(42, 8)),
	6497 => std_logic_vector(to_unsigned(42, 8)),
	6498 => std_logic_vector(to_unsigned(41, 8)),
	6499 => std_logic_vector(to_unsigned(41, 8)),
	6500 => std_logic_vector(to_unsigned(42, 8)),
	6501 => std_logic_vector(to_unsigned(41, 8)),
	6502 => std_logic_vector(to_unsigned(42, 8)),
	6503 => std_logic_vector(to_unsigned(42, 8)),
	6504 => std_logic_vector(to_unsigned(42, 8)),
	6505 => std_logic_vector(to_unsigned(42, 8)),
	6506 => std_logic_vector(to_unsigned(41, 8)),
	6507 => std_logic_vector(to_unsigned(42, 8)),
	6508 => std_logic_vector(to_unsigned(42, 8)),
	6509 => std_logic_vector(to_unsigned(42, 8)),
	6510 => std_logic_vector(to_unsigned(42, 8)),
	6511 => std_logic_vector(to_unsigned(41, 8)),
	6512 => std_logic_vector(to_unsigned(41, 8)),
	6513 => std_logic_vector(to_unsigned(42, 8)),
	6514 => std_logic_vector(to_unsigned(41, 8)),
	6515 => std_logic_vector(to_unsigned(42, 8)),
	6516 => std_logic_vector(to_unsigned(42, 8)),
	6517 => std_logic_vector(to_unsigned(41, 8)),
	6518 => std_logic_vector(to_unsigned(41, 8)),
	6519 => std_logic_vector(to_unsigned(41, 8)),
	6520 => std_logic_vector(to_unsigned(42, 8)),
	6521 => std_logic_vector(to_unsigned(42, 8)),
	6522 => std_logic_vector(to_unsigned(41, 8)),
	6523 => std_logic_vector(to_unsigned(42, 8)),
	6524 => std_logic_vector(to_unsigned(42, 8)),
	6525 => std_logic_vector(to_unsigned(41, 8)),
	6526 => std_logic_vector(to_unsigned(41, 8)),
	6527 => std_logic_vector(to_unsigned(41, 8)),
	6528 => std_logic_vector(to_unsigned(41, 8)),
	6529 => std_logic_vector(to_unsigned(42, 8)),
	6530 => std_logic_vector(to_unsigned(42, 8)),
	6531 => std_logic_vector(to_unsigned(42, 8)),
	6532 => std_logic_vector(to_unsigned(41, 8)),
	6533 => std_logic_vector(to_unsigned(41, 8)),
	6534 => std_logic_vector(to_unsigned(41, 8)),
	6535 => std_logic_vector(to_unsigned(41, 8)),
	6536 => std_logic_vector(to_unsigned(41, 8)),
	6537 => std_logic_vector(to_unsigned(41, 8)),
	6538 => std_logic_vector(to_unsigned(42, 8)),
	6539 => std_logic_vector(to_unsigned(42, 8)),
	6540 => std_logic_vector(to_unsigned(41, 8)),
	6541 => std_logic_vector(to_unsigned(41, 8)),
	6542 => std_logic_vector(to_unsigned(42, 8)),
	6543 => std_logic_vector(to_unsigned(41, 8)),
	6544 => std_logic_vector(to_unsigned(41, 8)),
	6545 => std_logic_vector(to_unsigned(42, 8)),
	6546 => std_logic_vector(to_unsigned(42, 8)),
	6547 => std_logic_vector(to_unsigned(42, 8)),
	6548 => std_logic_vector(to_unsigned(42, 8)),
	6549 => std_logic_vector(to_unsigned(42, 8)),
	6550 => std_logic_vector(to_unsigned(42, 8)),
	6551 => std_logic_vector(to_unsigned(42, 8)),
	6552 => std_logic_vector(to_unsigned(41, 8)),
	6553 => std_logic_vector(to_unsigned(42, 8)),
	6554 => std_logic_vector(to_unsigned(41, 8)),
	6555 => std_logic_vector(to_unsigned(42, 8)),
	6556 => std_logic_vector(to_unsigned(42, 8)),
	6557 => std_logic_vector(to_unsigned(41, 8)),
	6558 => std_logic_vector(to_unsigned(42, 8)),
	6559 => std_logic_vector(to_unsigned(42, 8)),
	6560 => std_logic_vector(to_unsigned(42, 8)),
	6561 => std_logic_vector(to_unsigned(42, 8)),
	6562 => std_logic_vector(to_unsigned(41, 8)),
	6563 => std_logic_vector(to_unsigned(42, 8)),
	6564 => std_logic_vector(to_unsigned(41, 8)),
	6565 => std_logic_vector(to_unsigned(42, 8)),
	6566 => std_logic_vector(to_unsigned(42, 8)),
	6567 => std_logic_vector(to_unsigned(41, 8)),
	6568 => std_logic_vector(to_unsigned(41, 8)),
	6569 => std_logic_vector(to_unsigned(41, 8)),
	6570 => std_logic_vector(to_unsigned(42, 8)),
	6571 => std_logic_vector(to_unsigned(42, 8)),
	6572 => std_logic_vector(to_unsigned(42, 8)),
	6573 => std_logic_vector(to_unsigned(41, 8)),
	6574 => std_logic_vector(to_unsigned(42, 8)),
	6575 => std_logic_vector(to_unsigned(42, 8)),
	6576 => std_logic_vector(to_unsigned(42, 8)),
	6577 => std_logic_vector(to_unsigned(42, 8)),
	6578 => std_logic_vector(to_unsigned(41, 8)),
	6579 => std_logic_vector(to_unsigned(41, 8)),
	6580 => std_logic_vector(to_unsigned(42, 8)),
	6581 => std_logic_vector(to_unsigned(42, 8)),
	6582 => std_logic_vector(to_unsigned(42, 8)),
	6583 => std_logic_vector(to_unsigned(42, 8)),
	6584 => std_logic_vector(to_unsigned(42, 8)),
	6585 => std_logic_vector(to_unsigned(42, 8)),
	6586 => std_logic_vector(to_unsigned(41, 8)),
	6587 => std_logic_vector(to_unsigned(42, 8)),
	6588 => std_logic_vector(to_unsigned(42, 8)),
	6589 => std_logic_vector(to_unsigned(42, 8)),
	6590 => std_logic_vector(to_unsigned(41, 8)),
	6591 => std_logic_vector(to_unsigned(42, 8)),
	6592 => std_logic_vector(to_unsigned(42, 8)),
	6593 => std_logic_vector(to_unsigned(41, 8)),
	6594 => std_logic_vector(to_unsigned(41, 8)),
	6595 => std_logic_vector(to_unsigned(42, 8)),
	6596 => std_logic_vector(to_unsigned(42, 8)),
	6597 => std_logic_vector(to_unsigned(41, 8)),
	6598 => std_logic_vector(to_unsigned(42, 8)),
	6599 => std_logic_vector(to_unsigned(42, 8)),
	6600 => std_logic_vector(to_unsigned(42, 8)),
	6601 => std_logic_vector(to_unsigned(41, 8)),
	6602 => std_logic_vector(to_unsigned(41, 8)),
	6603 => std_logic_vector(to_unsigned(41, 8)),
	6604 => std_logic_vector(to_unsigned(41, 8)),
	6605 => std_logic_vector(to_unsigned(41, 8)),
	6606 => std_logic_vector(to_unsigned(42, 8)),
	6607 => std_logic_vector(to_unsigned(42, 8)),
	6608 => std_logic_vector(to_unsigned(42, 8)),
	6609 => std_logic_vector(to_unsigned(41, 8)),
	6610 => std_logic_vector(to_unsigned(41, 8)),
	6611 => std_logic_vector(to_unsigned(42, 8)),
	6612 => std_logic_vector(to_unsigned(41, 8)),
	6613 => std_logic_vector(to_unsigned(42, 8)),
	6614 => std_logic_vector(to_unsigned(41, 8)),
	6615 => std_logic_vector(to_unsigned(41, 8)),
	6616 => std_logic_vector(to_unsigned(42, 8)),
	6617 => std_logic_vector(to_unsigned(42, 8)),
	6618 => std_logic_vector(to_unsigned(41, 8)),
	6619 => std_logic_vector(to_unsigned(42, 8)),
	6620 => std_logic_vector(to_unsigned(41, 8)),
	6621 => std_logic_vector(to_unsigned(42, 8)),
	6622 => std_logic_vector(to_unsigned(41, 8)),
	6623 => std_logic_vector(to_unsigned(42, 8)),
	6624 => std_logic_vector(to_unsigned(41, 8)),
	6625 => std_logic_vector(to_unsigned(41, 8)),
	6626 => std_logic_vector(to_unsigned(41, 8)),
	6627 => std_logic_vector(to_unsigned(42, 8)),
	6628 => std_logic_vector(to_unsigned(42, 8)),
	6629 => std_logic_vector(to_unsigned(42, 8)),
	6630 => std_logic_vector(to_unsigned(42, 8)),
	6631 => std_logic_vector(to_unsigned(42, 8)),
	6632 => std_logic_vector(to_unsigned(41, 8)),
	6633 => std_logic_vector(to_unsigned(42, 8)),
	6634 => std_logic_vector(to_unsigned(42, 8)),
	6635 => std_logic_vector(to_unsigned(42, 8)),
	6636 => std_logic_vector(to_unsigned(41, 8)),
	6637 => std_logic_vector(to_unsigned(42, 8)),
	6638 => std_logic_vector(to_unsigned(42, 8)),
	6639 => std_logic_vector(to_unsigned(41, 8)),
	6640 => std_logic_vector(to_unsigned(42, 8)),
	6641 => std_logic_vector(to_unsigned(41, 8)),
	6642 => std_logic_vector(to_unsigned(41, 8)),
	6643 => std_logic_vector(to_unsigned(41, 8)),
	6644 => std_logic_vector(to_unsigned(42, 8)),
	6645 => std_logic_vector(to_unsigned(42, 8)),
	6646 => std_logic_vector(to_unsigned(42, 8)),
	6647 => std_logic_vector(to_unsigned(41, 8)),
	6648 => std_logic_vector(to_unsigned(41, 8)),
	6649 => std_logic_vector(to_unsigned(41, 8)),
	6650 => std_logic_vector(to_unsigned(41, 8)),
	6651 => std_logic_vector(to_unsigned(41, 8)),
	6652 => std_logic_vector(to_unsigned(41, 8)),
	6653 => std_logic_vector(to_unsigned(42, 8)),
	6654 => std_logic_vector(to_unsigned(41, 8)),
	6655 => std_logic_vector(to_unsigned(41, 8)),
	6656 => std_logic_vector(to_unsigned(42, 8)),
	6657 => std_logic_vector(to_unsigned(41, 8)),
	6658 => std_logic_vector(to_unsigned(41, 8)),
	6659 => std_logic_vector(to_unsigned(42, 8)),
	6660 => std_logic_vector(to_unsigned(42, 8)),
	6661 => std_logic_vector(to_unsigned(41, 8)),
	6662 => std_logic_vector(to_unsigned(41, 8)),
	6663 => std_logic_vector(to_unsigned(41, 8)),
	6664 => std_logic_vector(to_unsigned(42, 8)),
	6665 => std_logic_vector(to_unsigned(42, 8)),
	6666 => std_logic_vector(to_unsigned(42, 8)),
	6667 => std_logic_vector(to_unsigned(42, 8)),
	6668 => std_logic_vector(to_unsigned(42, 8)),
	6669 => std_logic_vector(to_unsigned(41, 8)),
	6670 => std_logic_vector(to_unsigned(42, 8)),
	6671 => std_logic_vector(to_unsigned(41, 8)),
	6672 => std_logic_vector(to_unsigned(41, 8)),
	6673 => std_logic_vector(to_unsigned(42, 8)),
	6674 => std_logic_vector(to_unsigned(42, 8)),
	6675 => std_logic_vector(to_unsigned(41, 8)),
	6676 => std_logic_vector(to_unsigned(41, 8)),
	6677 => std_logic_vector(to_unsigned(42, 8)),
	6678 => std_logic_vector(to_unsigned(41, 8)),
	6679 => std_logic_vector(to_unsigned(42, 8)),
	6680 => std_logic_vector(to_unsigned(42, 8)),
	6681 => std_logic_vector(to_unsigned(42, 8)),
	6682 => std_logic_vector(to_unsigned(42, 8)),
	6683 => std_logic_vector(to_unsigned(41, 8)),
	6684 => std_logic_vector(to_unsigned(41, 8)),
	6685 => std_logic_vector(to_unsigned(42, 8)),
	6686 => std_logic_vector(to_unsigned(41, 8)),
	6687 => std_logic_vector(to_unsigned(41, 8)),
	6688 => std_logic_vector(to_unsigned(42, 8)),
	6689 => std_logic_vector(to_unsigned(41, 8)),
	6690 => std_logic_vector(to_unsigned(42, 8)),
	6691 => std_logic_vector(to_unsigned(41, 8)),
	6692 => std_logic_vector(to_unsigned(42, 8)),
	6693 => std_logic_vector(to_unsigned(41, 8)),
	6694 => std_logic_vector(to_unsigned(41, 8)),
	6695 => std_logic_vector(to_unsigned(41, 8)),
	6696 => std_logic_vector(to_unsigned(42, 8)),
	6697 => std_logic_vector(to_unsigned(41, 8)),
	6698 => std_logic_vector(to_unsigned(41, 8)),
	6699 => std_logic_vector(to_unsigned(42, 8)),
	6700 => std_logic_vector(to_unsigned(42, 8)),
	6701 => std_logic_vector(to_unsigned(41, 8)),
	6702 => std_logic_vector(to_unsigned(42, 8)),
	6703 => std_logic_vector(to_unsigned(41, 8)),
	6704 => std_logic_vector(to_unsigned(41, 8)),
	6705 => std_logic_vector(to_unsigned(42, 8)),
	6706 => std_logic_vector(to_unsigned(42, 8)),
	6707 => std_logic_vector(to_unsigned(42, 8)),
	6708 => std_logic_vector(to_unsigned(42, 8)),
	6709 => std_logic_vector(to_unsigned(41, 8)),
	6710 => std_logic_vector(to_unsigned(41, 8)),
	6711 => std_logic_vector(to_unsigned(41, 8)),
	6712 => std_logic_vector(to_unsigned(41, 8)),
	6713 => std_logic_vector(to_unsigned(42, 8)),
	6714 => std_logic_vector(to_unsigned(42, 8)),
	6715 => std_logic_vector(to_unsigned(41, 8)),
	6716 => std_logic_vector(to_unsigned(41, 8)),
	6717 => std_logic_vector(to_unsigned(41, 8)),
	others =>(others =>'0'));

component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_rst         : in  std_logic;
      i_start       : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector (7 downto 0)
      );
end component project_reti_logiche;


begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_rst      	=> tb_rst,
          i_start       => tb_start,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
          o_we 		=> mem_we,
          o_data    	=> mem_i_data
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;


MEM : process(tb_clk)
begin
    if tb_clk'event and tb_clk = '1' then
        if enable_wire = '1' then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
            end if;
        end if;
    end if;
end process;


test : process is
begin
    wait for 100 ns;
    wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_rst <= '0';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;

    assert RAM(6718) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6718)))) severity failure;
    assert RAM(6719) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6719)))) severity failure;
    assert RAM(6720) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6720)))) severity failure;
    assert RAM(6721) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6721)))) severity failure;
    assert RAM(6722) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6722)))) severity failure;
    assert RAM(6723) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6723)))) severity failure;
    assert RAM(6724) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6724)))) severity failure;
    assert RAM(6725) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6725)))) severity failure;
    assert RAM(6726) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6726)))) severity failure;
    assert RAM(6727) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6727)))) severity failure;
    assert RAM(6728) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6728)))) severity failure;
    assert RAM(6729) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6729)))) severity failure;
    assert RAM(6730) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6730)))) severity failure;
    assert RAM(6731) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6731)))) severity failure;
    assert RAM(6732) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6732)))) severity failure;
    assert RAM(6733) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6733)))) severity failure;
    assert RAM(6734) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6734)))) severity failure;
    assert RAM(6735) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6735)))) severity failure;
    assert RAM(6736) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6736)))) severity failure;
    assert RAM(6737) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6737)))) severity failure;
    assert RAM(6738) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6738)))) severity failure;
    assert RAM(6739) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6739)))) severity failure;
    assert RAM(6740) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6740)))) severity failure;
    assert RAM(6741) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6741)))) severity failure;
    assert RAM(6742) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6742)))) severity failure;
    assert RAM(6743) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6743)))) severity failure;
    assert RAM(6744) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6744)))) severity failure;
    assert RAM(6745) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6745)))) severity failure;
    assert RAM(6746) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6746)))) severity failure;
    assert RAM(6747) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6747)))) severity failure;
    assert RAM(6748) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6748)))) severity failure;
    assert RAM(6749) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6749)))) severity failure;
    assert RAM(6750) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6750)))) severity failure;
    assert RAM(6751) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6751)))) severity failure;
    assert RAM(6752) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6752)))) severity failure;
    assert RAM(6753) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6753)))) severity failure;
    assert RAM(6754) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6754)))) severity failure;
    assert RAM(6755) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6755)))) severity failure;
    assert RAM(6756) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6756)))) severity failure;
    assert RAM(6757) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6757)))) severity failure;
    assert RAM(6758) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6758)))) severity failure;
    assert RAM(6759) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6759)))) severity failure;
    assert RAM(6760) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6760)))) severity failure;
    assert RAM(6761) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6761)))) severity failure;
    assert RAM(6762) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6762)))) severity failure;
    assert RAM(6763) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6763)))) severity failure;
    assert RAM(6764) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6764)))) severity failure;
    assert RAM(6765) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6765)))) severity failure;
    assert RAM(6766) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6766)))) severity failure;
    assert RAM(6767) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6767)))) severity failure;
    assert RAM(6768) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6768)))) severity failure;
    assert RAM(6769) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6769)))) severity failure;
    assert RAM(6770) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6770)))) severity failure;
    assert RAM(6771) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6771)))) severity failure;
    assert RAM(6772) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6772)))) severity failure;
    assert RAM(6773) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6773)))) severity failure;
    assert RAM(6774) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6774)))) severity failure;
    assert RAM(6775) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6775)))) severity failure;
    assert RAM(6776) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6776)))) severity failure;
    assert RAM(6777) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6777)))) severity failure;
    assert RAM(6778) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6778)))) severity failure;
    assert RAM(6779) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6779)))) severity failure;
    assert RAM(6780) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6780)))) severity failure;
    assert RAM(6781) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6781)))) severity failure;
    assert RAM(6782) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6782)))) severity failure;
    assert RAM(6783) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6783)))) severity failure;
    assert RAM(6784) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6784)))) severity failure;
    assert RAM(6785) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6785)))) severity failure;
    assert RAM(6786) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6786)))) severity failure;
    assert RAM(6787) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6787)))) severity failure;
    assert RAM(6788) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6788)))) severity failure;
    assert RAM(6789) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6789)))) severity failure;
    assert RAM(6790) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6790)))) severity failure;
    assert RAM(6791) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6791)))) severity failure;
    assert RAM(6792) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6792)))) severity failure;
    assert RAM(6793) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6793)))) severity failure;
    assert RAM(6794) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6794)))) severity failure;
    assert RAM(6795) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6795)))) severity failure;
    assert RAM(6796) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6796)))) severity failure;
    assert RAM(6797) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6797)))) severity failure;
    assert RAM(6798) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6798)))) severity failure;
    assert RAM(6799) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6799)))) severity failure;
    assert RAM(6800) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6800)))) severity failure;
    assert RAM(6801) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6801)))) severity failure;
    assert RAM(6802) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6802)))) severity failure;
    assert RAM(6803) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6803)))) severity failure;
    assert RAM(6804) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6804)))) severity failure;
    assert RAM(6805) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6805)))) severity failure;
    assert RAM(6806) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6806)))) severity failure;
    assert RAM(6807) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6807)))) severity failure;
    assert RAM(6808) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6808)))) severity failure;
    assert RAM(6809) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6809)))) severity failure;
    assert RAM(6810) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6810)))) severity failure;
    assert RAM(6811) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6811)))) severity failure;
    assert RAM(6812) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6812)))) severity failure;
    assert RAM(6813) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6813)))) severity failure;
    assert RAM(6814) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6814)))) severity failure;
    assert RAM(6815) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6815)))) severity failure;
    assert RAM(6816) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6816)))) severity failure;
    assert RAM(6817) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6817)))) severity failure;
    assert RAM(6818) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6818)))) severity failure;
    assert RAM(6819) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6819)))) severity failure;
    assert RAM(6820) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6820)))) severity failure;
    assert RAM(6821) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6821)))) severity failure;
    assert RAM(6822) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6822)))) severity failure;
    assert RAM(6823) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6823)))) severity failure;
    assert RAM(6824) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6824)))) severity failure;
    assert RAM(6825) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6825)))) severity failure;
    assert RAM(6826) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6826)))) severity failure;
    assert RAM(6827) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6827)))) severity failure;
    assert RAM(6828) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6828)))) severity failure;
    assert RAM(6829) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6829)))) severity failure;
    assert RAM(6830) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6830)))) severity failure;
    assert RAM(6831) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6831)))) severity failure;
    assert RAM(6832) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6832)))) severity failure;
    assert RAM(6833) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6833)))) severity failure;
    assert RAM(6834) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6834)))) severity failure;
    assert RAM(6835) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6835)))) severity failure;
    assert RAM(6836) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6836)))) severity failure;
    assert RAM(6837) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6837)))) severity failure;
    assert RAM(6838) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6838)))) severity failure;
    assert RAM(6839) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6839)))) severity failure;
    assert RAM(6840) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6840)))) severity failure;
    assert RAM(6841) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6841)))) severity failure;
    assert RAM(6842) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6842)))) severity failure;
    assert RAM(6843) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6843)))) severity failure;
    assert RAM(6844) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6844)))) severity failure;
    assert RAM(6845) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6845)))) severity failure;
    assert RAM(6846) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6846)))) severity failure;
    assert RAM(6847) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6847)))) severity failure;
    assert RAM(6848) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6848)))) severity failure;
    assert RAM(6849) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6849)))) severity failure;
    assert RAM(6850) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6850)))) severity failure;
    assert RAM(6851) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6851)))) severity failure;
    assert RAM(6852) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6852)))) severity failure;
    assert RAM(6853) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6853)))) severity failure;
    assert RAM(6854) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6854)))) severity failure;
    assert RAM(6855) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6855)))) severity failure;
    assert RAM(6856) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6856)))) severity failure;
    assert RAM(6857) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6857)))) severity failure;
    assert RAM(6858) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6858)))) severity failure;
    assert RAM(6859) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6859)))) severity failure;
    assert RAM(6860) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6860)))) severity failure;
    assert RAM(6861) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6861)))) severity failure;
    assert RAM(6862) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6862)))) severity failure;
    assert RAM(6863) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6863)))) severity failure;
    assert RAM(6864) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6864)))) severity failure;
    assert RAM(6865) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6865)))) severity failure;
    assert RAM(6866) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6866)))) severity failure;
    assert RAM(6867) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6867)))) severity failure;
    assert RAM(6868) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6868)))) severity failure;
    assert RAM(6869) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6869)))) severity failure;
    assert RAM(6870) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6870)))) severity failure;
    assert RAM(6871) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6871)))) severity failure;
    assert RAM(6872) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6872)))) severity failure;
    assert RAM(6873) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6873)))) severity failure;
    assert RAM(6874) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6874)))) severity failure;
    assert RAM(6875) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6875)))) severity failure;
    assert RAM(6876) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6876)))) severity failure;
    assert RAM(6877) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6877)))) severity failure;
    assert RAM(6878) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6878)))) severity failure;
    assert RAM(6879) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6879)))) severity failure;
    assert RAM(6880) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6880)))) severity failure;
    assert RAM(6881) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6881)))) severity failure;
    assert RAM(6882) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6882)))) severity failure;
    assert RAM(6883) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6883)))) severity failure;
    assert RAM(6884) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6884)))) severity failure;
    assert RAM(6885) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6885)))) severity failure;
    assert RAM(6886) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6886)))) severity failure;
    assert RAM(6887) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6887)))) severity failure;
    assert RAM(6888) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6888)))) severity failure;
    assert RAM(6889) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6889)))) severity failure;
    assert RAM(6890) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6890)))) severity failure;
    assert RAM(6891) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6891)))) severity failure;
    assert RAM(6892) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6892)))) severity failure;
    assert RAM(6893) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6893)))) severity failure;
    assert RAM(6894) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6894)))) severity failure;
    assert RAM(6895) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6895)))) severity failure;
    assert RAM(6896) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6896)))) severity failure;
    assert RAM(6897) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6897)))) severity failure;
    assert RAM(6898) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6898)))) severity failure;
    assert RAM(6899) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6899)))) severity failure;
    assert RAM(6900) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6900)))) severity failure;
    assert RAM(6901) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6901)))) severity failure;
    assert RAM(6902) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6902)))) severity failure;
    assert RAM(6903) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6903)))) severity failure;
    assert RAM(6904) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6904)))) severity failure;
    assert RAM(6905) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6905)))) severity failure;
    assert RAM(6906) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6906)))) severity failure;
    assert RAM(6907) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6907)))) severity failure;
    assert RAM(6908) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6908)))) severity failure;
    assert RAM(6909) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6909)))) severity failure;
    assert RAM(6910) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6910)))) severity failure;
    assert RAM(6911) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6911)))) severity failure;
    assert RAM(6912) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6912)))) severity failure;
    assert RAM(6913) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6913)))) severity failure;
    assert RAM(6914) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6914)))) severity failure;
    assert RAM(6915) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6915)))) severity failure;
    assert RAM(6916) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6916)))) severity failure;
    assert RAM(6917) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6917)))) severity failure;
    assert RAM(6918) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6918)))) severity failure;
    assert RAM(6919) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6919)))) severity failure;
    assert RAM(6920) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6920)))) severity failure;
    assert RAM(6921) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6921)))) severity failure;
    assert RAM(6922) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6922)))) severity failure;
    assert RAM(6923) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6923)))) severity failure;
    assert RAM(6924) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6924)))) severity failure;
    assert RAM(6925) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6925)))) severity failure;
    assert RAM(6926) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6926)))) severity failure;
    assert RAM(6927) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6927)))) severity failure;
    assert RAM(6928) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6928)))) severity failure;
    assert RAM(6929) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6929)))) severity failure;
    assert RAM(6930) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6930)))) severity failure;
    assert RAM(6931) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6931)))) severity failure;
    assert RAM(6932) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6932)))) severity failure;
    assert RAM(6933) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6933)))) severity failure;
    assert RAM(6934) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6934)))) severity failure;
    assert RAM(6935) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6935)))) severity failure;
    assert RAM(6936) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6936)))) severity failure;
    assert RAM(6937) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6937)))) severity failure;
    assert RAM(6938) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6938)))) severity failure;
    assert RAM(6939) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6939)))) severity failure;
    assert RAM(6940) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6940)))) severity failure;
    assert RAM(6941) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6941)))) severity failure;
    assert RAM(6942) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6942)))) severity failure;
    assert RAM(6943) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6943)))) severity failure;
    assert RAM(6944) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6944)))) severity failure;
    assert RAM(6945) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6945)))) severity failure;
    assert RAM(6946) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6946)))) severity failure;
    assert RAM(6947) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6947)))) severity failure;
    assert RAM(6948) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6948)))) severity failure;
    assert RAM(6949) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6949)))) severity failure;
    assert RAM(6950) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6950)))) severity failure;
    assert RAM(6951) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6951)))) severity failure;
    assert RAM(6952) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6952)))) severity failure;
    assert RAM(6953) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6953)))) severity failure;
    assert RAM(6954) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6954)))) severity failure;
    assert RAM(6955) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6955)))) severity failure;
    assert RAM(6956) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6956)))) severity failure;
    assert RAM(6957) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6957)))) severity failure;
    assert RAM(6958) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6958)))) severity failure;
    assert RAM(6959) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6959)))) severity failure;
    assert RAM(6960) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6960)))) severity failure;
    assert RAM(6961) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6961)))) severity failure;
    assert RAM(6962) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6962)))) severity failure;
    assert RAM(6963) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6963)))) severity failure;
    assert RAM(6964) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6964)))) severity failure;
    assert RAM(6965) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6965)))) severity failure;
    assert RAM(6966) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6966)))) severity failure;
    assert RAM(6967) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6967)))) severity failure;
    assert RAM(6968) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6968)))) severity failure;
    assert RAM(6969) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6969)))) severity failure;
    assert RAM(6970) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6970)))) severity failure;
    assert RAM(6971) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6971)))) severity failure;
    assert RAM(6972) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6972)))) severity failure;
    assert RAM(6973) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6973)))) severity failure;
    assert RAM(6974) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6974)))) severity failure;
    assert RAM(6975) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6975)))) severity failure;
    assert RAM(6976) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6976)))) severity failure;
    assert RAM(6977) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6977)))) severity failure;
    assert RAM(6978) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6978)))) severity failure;
    assert RAM(6979) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6979)))) severity failure;
    assert RAM(6980) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6980)))) severity failure;
    assert RAM(6981) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6981)))) severity failure;
    assert RAM(6982) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6982)))) severity failure;
    assert RAM(6983) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6983)))) severity failure;
    assert RAM(6984) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6984)))) severity failure;
    assert RAM(6985) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6985)))) severity failure;
    assert RAM(6986) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6986)))) severity failure;
    assert RAM(6987) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6987)))) severity failure;
    assert RAM(6988) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6988)))) severity failure;
    assert RAM(6989) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6989)))) severity failure;
    assert RAM(6990) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6990)))) severity failure;
    assert RAM(6991) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6991)))) severity failure;
    assert RAM(6992) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(6992)))) severity failure;
    assert RAM(6993) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6993)))) severity failure;
    assert RAM(6994) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6994)))) severity failure;
    assert RAM(6995) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6995)))) severity failure;
    assert RAM(6996) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6996)))) severity failure;
    assert RAM(6997) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6997)))) severity failure;
    assert RAM(6998) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6998)))) severity failure;
    assert RAM(6999) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(6999)))) severity failure;
    assert RAM(7000) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7000)))) severity failure;
    assert RAM(7001) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7001)))) severity failure;
    assert RAM(7002) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7002)))) severity failure;
    assert RAM(7003) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7003)))) severity failure;
    assert RAM(7004) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7004)))) severity failure;
    assert RAM(7005) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7005)))) severity failure;
    assert RAM(7006) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7006)))) severity failure;
    assert RAM(7007) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7007)))) severity failure;
    assert RAM(7008) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7008)))) severity failure;
    assert RAM(7009) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7009)))) severity failure;
    assert RAM(7010) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7010)))) severity failure;
    assert RAM(7011) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7011)))) severity failure;
    assert RAM(7012) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7012)))) severity failure;
    assert RAM(7013) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7013)))) severity failure;
    assert RAM(7014) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7014)))) severity failure;
    assert RAM(7015) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7015)))) severity failure;
    assert RAM(7016) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7016)))) severity failure;
    assert RAM(7017) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7017)))) severity failure;
    assert RAM(7018) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7018)))) severity failure;
    assert RAM(7019) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7019)))) severity failure;
    assert RAM(7020) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7020)))) severity failure;
    assert RAM(7021) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7021)))) severity failure;
    assert RAM(7022) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7022)))) severity failure;
    assert RAM(7023) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7023)))) severity failure;
    assert RAM(7024) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7024)))) severity failure;
    assert RAM(7025) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7025)))) severity failure;
    assert RAM(7026) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7026)))) severity failure;
    assert RAM(7027) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7027)))) severity failure;
    assert RAM(7028) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7028)))) severity failure;
    assert RAM(7029) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7029)))) severity failure;
    assert RAM(7030) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7030)))) severity failure;
    assert RAM(7031) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7031)))) severity failure;
    assert RAM(7032) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7032)))) severity failure;
    assert RAM(7033) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7033)))) severity failure;
    assert RAM(7034) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7034)))) severity failure;
    assert RAM(7035) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7035)))) severity failure;
    assert RAM(7036) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7036)))) severity failure;
    assert RAM(7037) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7037)))) severity failure;
    assert RAM(7038) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7038)))) severity failure;
    assert RAM(7039) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7039)))) severity failure;
    assert RAM(7040) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7040)))) severity failure;
    assert RAM(7041) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7041)))) severity failure;
    assert RAM(7042) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7042)))) severity failure;
    assert RAM(7043) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7043)))) severity failure;
    assert RAM(7044) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7044)))) severity failure;
    assert RAM(7045) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7045)))) severity failure;
    assert RAM(7046) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7046)))) severity failure;
    assert RAM(7047) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7047)))) severity failure;
    assert RAM(7048) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7048)))) severity failure;
    assert RAM(7049) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7049)))) severity failure;
    assert RAM(7050) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7050)))) severity failure;
    assert RAM(7051) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7051)))) severity failure;
    assert RAM(7052) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7052)))) severity failure;
    assert RAM(7053) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7053)))) severity failure;
    assert RAM(7054) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7054)))) severity failure;
    assert RAM(7055) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7055)))) severity failure;
    assert RAM(7056) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7056)))) severity failure;
    assert RAM(7057) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7057)))) severity failure;
    assert RAM(7058) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7058)))) severity failure;
    assert RAM(7059) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7059)))) severity failure;
    assert RAM(7060) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7060)))) severity failure;
    assert RAM(7061) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7061)))) severity failure;
    assert RAM(7062) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7062)))) severity failure;
    assert RAM(7063) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7063)))) severity failure;
    assert RAM(7064) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7064)))) severity failure;
    assert RAM(7065) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7065)))) severity failure;
    assert RAM(7066) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7066)))) severity failure;
    assert RAM(7067) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7067)))) severity failure;
    assert RAM(7068) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7068)))) severity failure;
    assert RAM(7069) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7069)))) severity failure;
    assert RAM(7070) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7070)))) severity failure;
    assert RAM(7071) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7071)))) severity failure;
    assert RAM(7072) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7072)))) severity failure;
    assert RAM(7073) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7073)))) severity failure;
    assert RAM(7074) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7074)))) severity failure;
    assert RAM(7075) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7075)))) severity failure;
    assert RAM(7076) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7076)))) severity failure;
    assert RAM(7077) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7077)))) severity failure;
    assert RAM(7078) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7078)))) severity failure;
    assert RAM(7079) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7079)))) severity failure;
    assert RAM(7080) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7080)))) severity failure;
    assert RAM(7081) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7081)))) severity failure;
    assert RAM(7082) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7082)))) severity failure;
    assert RAM(7083) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7083)))) severity failure;
    assert RAM(7084) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7084)))) severity failure;
    assert RAM(7085) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7085)))) severity failure;
    assert RAM(7086) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7086)))) severity failure;
    assert RAM(7087) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7087)))) severity failure;
    assert RAM(7088) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7088)))) severity failure;
    assert RAM(7089) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7089)))) severity failure;
    assert RAM(7090) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7090)))) severity failure;
    assert RAM(7091) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7091)))) severity failure;
    assert RAM(7092) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7092)))) severity failure;
    assert RAM(7093) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7093)))) severity failure;
    assert RAM(7094) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7094)))) severity failure;
    assert RAM(7095) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7095)))) severity failure;
    assert RAM(7096) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7096)))) severity failure;
    assert RAM(7097) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7097)))) severity failure;
    assert RAM(7098) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7098)))) severity failure;
    assert RAM(7099) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7099)))) severity failure;
    assert RAM(7100) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7100)))) severity failure;
    assert RAM(7101) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7101)))) severity failure;
    assert RAM(7102) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7102)))) severity failure;
    assert RAM(7103) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7103)))) severity failure;
    assert RAM(7104) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7104)))) severity failure;
    assert RAM(7105) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7105)))) severity failure;
    assert RAM(7106) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7106)))) severity failure;
    assert RAM(7107) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7107)))) severity failure;
    assert RAM(7108) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7108)))) severity failure;
    assert RAM(7109) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7109)))) severity failure;
    assert RAM(7110) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7110)))) severity failure;
    assert RAM(7111) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7111)))) severity failure;
    assert RAM(7112) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7112)))) severity failure;
    assert RAM(7113) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7113)))) severity failure;
    assert RAM(7114) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7114)))) severity failure;
    assert RAM(7115) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7115)))) severity failure;
    assert RAM(7116) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7116)))) severity failure;
    assert RAM(7117) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7117)))) severity failure;
    assert RAM(7118) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7118)))) severity failure;
    assert RAM(7119) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7119)))) severity failure;
    assert RAM(7120) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7120)))) severity failure;
    assert RAM(7121) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7121)))) severity failure;
    assert RAM(7122) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7122)))) severity failure;
    assert RAM(7123) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7123)))) severity failure;
    assert RAM(7124) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7124)))) severity failure;
    assert RAM(7125) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7125)))) severity failure;
    assert RAM(7126) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7126)))) severity failure;
    assert RAM(7127) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7127)))) severity failure;
    assert RAM(7128) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7128)))) severity failure;
    assert RAM(7129) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7129)))) severity failure;
    assert RAM(7130) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7130)))) severity failure;
    assert RAM(7131) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7131)))) severity failure;
    assert RAM(7132) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7132)))) severity failure;
    assert RAM(7133) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7133)))) severity failure;
    assert RAM(7134) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7134)))) severity failure;
    assert RAM(7135) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7135)))) severity failure;
    assert RAM(7136) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7136)))) severity failure;
    assert RAM(7137) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7137)))) severity failure;
    assert RAM(7138) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7138)))) severity failure;
    assert RAM(7139) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7139)))) severity failure;
    assert RAM(7140) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7140)))) severity failure;
    assert RAM(7141) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7141)))) severity failure;
    assert RAM(7142) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7142)))) severity failure;
    assert RAM(7143) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7143)))) severity failure;
    assert RAM(7144) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7144)))) severity failure;
    assert RAM(7145) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7145)))) severity failure;
    assert RAM(7146) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7146)))) severity failure;
    assert RAM(7147) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7147)))) severity failure;
    assert RAM(7148) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7148)))) severity failure;
    assert RAM(7149) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7149)))) severity failure;
    assert RAM(7150) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7150)))) severity failure;
    assert RAM(7151) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7151)))) severity failure;
    assert RAM(7152) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7152)))) severity failure;
    assert RAM(7153) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7153)))) severity failure;
    assert RAM(7154) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7154)))) severity failure;
    assert RAM(7155) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7155)))) severity failure;
    assert RAM(7156) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7156)))) severity failure;
    assert RAM(7157) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7157)))) severity failure;
    assert RAM(7158) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7158)))) severity failure;
    assert RAM(7159) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7159)))) severity failure;
    assert RAM(7160) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7160)))) severity failure;
    assert RAM(7161) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7161)))) severity failure;
    assert RAM(7162) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7162)))) severity failure;
    assert RAM(7163) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7163)))) severity failure;
    assert RAM(7164) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7164)))) severity failure;
    assert RAM(7165) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7165)))) severity failure;
    assert RAM(7166) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7166)))) severity failure;
    assert RAM(7167) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7167)))) severity failure;
    assert RAM(7168) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7168)))) severity failure;
    assert RAM(7169) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7169)))) severity failure;
    assert RAM(7170) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7170)))) severity failure;
    assert RAM(7171) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7171)))) severity failure;
    assert RAM(7172) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7172)))) severity failure;
    assert RAM(7173) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7173)))) severity failure;
    assert RAM(7174) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7174)))) severity failure;
    assert RAM(7175) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7175)))) severity failure;
    assert RAM(7176) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7176)))) severity failure;
    assert RAM(7177) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7177)))) severity failure;
    assert RAM(7178) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7178)))) severity failure;
    assert RAM(7179) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7179)))) severity failure;
    assert RAM(7180) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7180)))) severity failure;
    assert RAM(7181) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7181)))) severity failure;
    assert RAM(7182) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7182)))) severity failure;
    assert RAM(7183) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7183)))) severity failure;
    assert RAM(7184) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7184)))) severity failure;
    assert RAM(7185) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7185)))) severity failure;
    assert RAM(7186) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7186)))) severity failure;
    assert RAM(7187) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7187)))) severity failure;
    assert RAM(7188) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7188)))) severity failure;
    assert RAM(7189) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7189)))) severity failure;
    assert RAM(7190) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7190)))) severity failure;
    assert RAM(7191) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7191)))) severity failure;
    assert RAM(7192) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7192)))) severity failure;
    assert RAM(7193) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7193)))) severity failure;
    assert RAM(7194) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7194)))) severity failure;
    assert RAM(7195) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7195)))) severity failure;
    assert RAM(7196) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7196)))) severity failure;
    assert RAM(7197) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7197)))) severity failure;
    assert RAM(7198) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7198)))) severity failure;
    assert RAM(7199) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7199)))) severity failure;
    assert RAM(7200) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7200)))) severity failure;
    assert RAM(7201) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7201)))) severity failure;
    assert RAM(7202) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7202)))) severity failure;
    assert RAM(7203) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7203)))) severity failure;
    assert RAM(7204) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7204)))) severity failure;
    assert RAM(7205) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7205)))) severity failure;
    assert RAM(7206) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7206)))) severity failure;
    assert RAM(7207) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7207)))) severity failure;
    assert RAM(7208) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7208)))) severity failure;
    assert RAM(7209) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7209)))) severity failure;
    assert RAM(7210) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7210)))) severity failure;
    assert RAM(7211) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7211)))) severity failure;
    assert RAM(7212) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7212)))) severity failure;
    assert RAM(7213) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7213)))) severity failure;
    assert RAM(7214) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7214)))) severity failure;
    assert RAM(7215) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7215)))) severity failure;
    assert RAM(7216) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7216)))) severity failure;
    assert RAM(7217) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7217)))) severity failure;
    assert RAM(7218) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7218)))) severity failure;
    assert RAM(7219) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7219)))) severity failure;
    assert RAM(7220) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7220)))) severity failure;
    assert RAM(7221) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7221)))) severity failure;
    assert RAM(7222) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7222)))) severity failure;
    assert RAM(7223) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7223)))) severity failure;
    assert RAM(7224) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7224)))) severity failure;
    assert RAM(7225) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7225)))) severity failure;
    assert RAM(7226) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7226)))) severity failure;
    assert RAM(7227) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7227)))) severity failure;
    assert RAM(7228) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7228)))) severity failure;
    assert RAM(7229) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7229)))) severity failure;
    assert RAM(7230) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7230)))) severity failure;
    assert RAM(7231) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7231)))) severity failure;
    assert RAM(7232) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7232)))) severity failure;
    assert RAM(7233) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7233)))) severity failure;
    assert RAM(7234) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7234)))) severity failure;
    assert RAM(7235) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7235)))) severity failure;
    assert RAM(7236) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7236)))) severity failure;
    assert RAM(7237) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7237)))) severity failure;
    assert RAM(7238) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7238)))) severity failure;
    assert RAM(7239) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7239)))) severity failure;
    assert RAM(7240) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7240)))) severity failure;
    assert RAM(7241) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7241)))) severity failure;
    assert RAM(7242) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7242)))) severity failure;
    assert RAM(7243) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7243)))) severity failure;
    assert RAM(7244) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7244)))) severity failure;
    assert RAM(7245) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7245)))) severity failure;
    assert RAM(7246) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7246)))) severity failure;
    assert RAM(7247) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7247)))) severity failure;
    assert RAM(7248) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7248)))) severity failure;
    assert RAM(7249) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7249)))) severity failure;
    assert RAM(7250) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7250)))) severity failure;
    assert RAM(7251) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7251)))) severity failure;
    assert RAM(7252) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7252)))) severity failure;
    assert RAM(7253) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7253)))) severity failure;
    assert RAM(7254) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7254)))) severity failure;
    assert RAM(7255) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7255)))) severity failure;
    assert RAM(7256) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7256)))) severity failure;
    assert RAM(7257) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7257)))) severity failure;
    assert RAM(7258) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7258)))) severity failure;
    assert RAM(7259) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7259)))) severity failure;
    assert RAM(7260) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7260)))) severity failure;
    assert RAM(7261) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7261)))) severity failure;
    assert RAM(7262) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7262)))) severity failure;
    assert RAM(7263) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7263)))) severity failure;
    assert RAM(7264) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7264)))) severity failure;
    assert RAM(7265) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7265)))) severity failure;
    assert RAM(7266) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7266)))) severity failure;
    assert RAM(7267) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7267)))) severity failure;
    assert RAM(7268) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7268)))) severity failure;
    assert RAM(7269) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7269)))) severity failure;
    assert RAM(7270) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7270)))) severity failure;
    assert RAM(7271) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7271)))) severity failure;
    assert RAM(7272) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7272)))) severity failure;
    assert RAM(7273) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7273)))) severity failure;
    assert RAM(7274) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7274)))) severity failure;
    assert RAM(7275) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7275)))) severity failure;
    assert RAM(7276) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7276)))) severity failure;
    assert RAM(7277) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7277)))) severity failure;
    assert RAM(7278) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7278)))) severity failure;
    assert RAM(7279) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7279)))) severity failure;
    assert RAM(7280) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7280)))) severity failure;
    assert RAM(7281) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7281)))) severity failure;
    assert RAM(7282) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7282)))) severity failure;
    assert RAM(7283) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7283)))) severity failure;
    assert RAM(7284) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7284)))) severity failure;
    assert RAM(7285) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7285)))) severity failure;
    assert RAM(7286) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7286)))) severity failure;
    assert RAM(7287) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7287)))) severity failure;
    assert RAM(7288) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7288)))) severity failure;
    assert RAM(7289) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7289)))) severity failure;
    assert RAM(7290) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7290)))) severity failure;
    assert RAM(7291) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7291)))) severity failure;
    assert RAM(7292) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7292)))) severity failure;
    assert RAM(7293) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7293)))) severity failure;
    assert RAM(7294) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7294)))) severity failure;
    assert RAM(7295) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7295)))) severity failure;
    assert RAM(7296) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7296)))) severity failure;
    assert RAM(7297) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7297)))) severity failure;
    assert RAM(7298) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7298)))) severity failure;
    assert RAM(7299) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7299)))) severity failure;
    assert RAM(7300) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7300)))) severity failure;
    assert RAM(7301) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7301)))) severity failure;
    assert RAM(7302) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7302)))) severity failure;
    assert RAM(7303) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7303)))) severity failure;
    assert RAM(7304) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7304)))) severity failure;
    assert RAM(7305) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7305)))) severity failure;
    assert RAM(7306) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7306)))) severity failure;
    assert RAM(7307) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7307)))) severity failure;
    assert RAM(7308) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7308)))) severity failure;
    assert RAM(7309) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7309)))) severity failure;
    assert RAM(7310) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7310)))) severity failure;
    assert RAM(7311) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7311)))) severity failure;
    assert RAM(7312) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7312)))) severity failure;
    assert RAM(7313) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7313)))) severity failure;
    assert RAM(7314) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7314)))) severity failure;
    assert RAM(7315) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7315)))) severity failure;
    assert RAM(7316) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7316)))) severity failure;
    assert RAM(7317) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7317)))) severity failure;
    assert RAM(7318) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7318)))) severity failure;
    assert RAM(7319) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7319)))) severity failure;
    assert RAM(7320) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7320)))) severity failure;
    assert RAM(7321) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7321)))) severity failure;
    assert RAM(7322) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7322)))) severity failure;
    assert RAM(7323) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7323)))) severity failure;
    assert RAM(7324) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7324)))) severity failure;
    assert RAM(7325) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7325)))) severity failure;
    assert RAM(7326) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7326)))) severity failure;
    assert RAM(7327) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7327)))) severity failure;
    assert RAM(7328) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7328)))) severity failure;
    assert RAM(7329) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7329)))) severity failure;
    assert RAM(7330) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7330)))) severity failure;
    assert RAM(7331) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7331)))) severity failure;
    assert RAM(7332) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7332)))) severity failure;
    assert RAM(7333) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7333)))) severity failure;
    assert RAM(7334) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7334)))) severity failure;
    assert RAM(7335) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7335)))) severity failure;
    assert RAM(7336) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7336)))) severity failure;
    assert RAM(7337) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7337)))) severity failure;
    assert RAM(7338) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7338)))) severity failure;
    assert RAM(7339) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7339)))) severity failure;
    assert RAM(7340) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7340)))) severity failure;
    assert RAM(7341) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7341)))) severity failure;
    assert RAM(7342) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7342)))) severity failure;
    assert RAM(7343) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7343)))) severity failure;
    assert RAM(7344) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7344)))) severity failure;
    assert RAM(7345) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7345)))) severity failure;
    assert RAM(7346) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7346)))) severity failure;
    assert RAM(7347) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7347)))) severity failure;
    assert RAM(7348) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7348)))) severity failure;
    assert RAM(7349) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7349)))) severity failure;
    assert RAM(7350) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7350)))) severity failure;
    assert RAM(7351) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7351)))) severity failure;
    assert RAM(7352) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7352)))) severity failure;
    assert RAM(7353) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7353)))) severity failure;
    assert RAM(7354) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7354)))) severity failure;
    assert RAM(7355) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7355)))) severity failure;
    assert RAM(7356) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7356)))) severity failure;
    assert RAM(7357) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7357)))) severity failure;
    assert RAM(7358) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7358)))) severity failure;
    assert RAM(7359) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7359)))) severity failure;
    assert RAM(7360) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7360)))) severity failure;
    assert RAM(7361) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7361)))) severity failure;
    assert RAM(7362) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7362)))) severity failure;
    assert RAM(7363) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7363)))) severity failure;
    assert RAM(7364) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7364)))) severity failure;
    assert RAM(7365) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7365)))) severity failure;
    assert RAM(7366) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7366)))) severity failure;
    assert RAM(7367) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7367)))) severity failure;
    assert RAM(7368) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7368)))) severity failure;
    assert RAM(7369) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7369)))) severity failure;
    assert RAM(7370) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7370)))) severity failure;
    assert RAM(7371) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7371)))) severity failure;
    assert RAM(7372) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7372)))) severity failure;
    assert RAM(7373) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7373)))) severity failure;
    assert RAM(7374) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7374)))) severity failure;
    assert RAM(7375) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7375)))) severity failure;
    assert RAM(7376) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7376)))) severity failure;
    assert RAM(7377) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7377)))) severity failure;
    assert RAM(7378) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7378)))) severity failure;
    assert RAM(7379) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7379)))) severity failure;
    assert RAM(7380) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7380)))) severity failure;
    assert RAM(7381) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7381)))) severity failure;
    assert RAM(7382) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7382)))) severity failure;
    assert RAM(7383) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7383)))) severity failure;
    assert RAM(7384) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7384)))) severity failure;
    assert RAM(7385) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7385)))) severity failure;
    assert RAM(7386) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7386)))) severity failure;
    assert RAM(7387) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7387)))) severity failure;
    assert RAM(7388) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7388)))) severity failure;
    assert RAM(7389) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7389)))) severity failure;
    assert RAM(7390) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7390)))) severity failure;
    assert RAM(7391) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7391)))) severity failure;
    assert RAM(7392) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7392)))) severity failure;
    assert RAM(7393) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7393)))) severity failure;
    assert RAM(7394) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7394)))) severity failure;
    assert RAM(7395) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7395)))) severity failure;
    assert RAM(7396) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7396)))) severity failure;
    assert RAM(7397) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7397)))) severity failure;
    assert RAM(7398) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7398)))) severity failure;
    assert RAM(7399) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7399)))) severity failure;
    assert RAM(7400) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7400)))) severity failure;
    assert RAM(7401) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7401)))) severity failure;
    assert RAM(7402) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7402)))) severity failure;
    assert RAM(7403) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7403)))) severity failure;
    assert RAM(7404) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7404)))) severity failure;
    assert RAM(7405) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7405)))) severity failure;
    assert RAM(7406) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7406)))) severity failure;
    assert RAM(7407) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7407)))) severity failure;
    assert RAM(7408) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7408)))) severity failure;
    assert RAM(7409) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7409)))) severity failure;
    assert RAM(7410) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7410)))) severity failure;
    assert RAM(7411) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7411)))) severity failure;
    assert RAM(7412) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7412)))) severity failure;
    assert RAM(7413) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7413)))) severity failure;
    assert RAM(7414) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7414)))) severity failure;
    assert RAM(7415) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7415)))) severity failure;
    assert RAM(7416) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7416)))) severity failure;
    assert RAM(7417) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7417)))) severity failure;
    assert RAM(7418) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7418)))) severity failure;
    assert RAM(7419) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7419)))) severity failure;
    assert RAM(7420) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7420)))) severity failure;
    assert RAM(7421) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7421)))) severity failure;
    assert RAM(7422) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7422)))) severity failure;
    assert RAM(7423) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7423)))) severity failure;
    assert RAM(7424) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7424)))) severity failure;
    assert RAM(7425) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7425)))) severity failure;
    assert RAM(7426) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7426)))) severity failure;
    assert RAM(7427) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7427)))) severity failure;
    assert RAM(7428) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7428)))) severity failure;
    assert RAM(7429) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7429)))) severity failure;
    assert RAM(7430) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7430)))) severity failure;
    assert RAM(7431) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7431)))) severity failure;
    assert RAM(7432) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7432)))) severity failure;
    assert RAM(7433) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7433)))) severity failure;
    assert RAM(7434) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7434)))) severity failure;
    assert RAM(7435) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7435)))) severity failure;
    assert RAM(7436) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7436)))) severity failure;
    assert RAM(7437) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7437)))) severity failure;
    assert RAM(7438) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7438)))) severity failure;
    assert RAM(7439) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7439)))) severity failure;
    assert RAM(7440) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7440)))) severity failure;
    assert RAM(7441) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7441)))) severity failure;
    assert RAM(7442) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7442)))) severity failure;
    assert RAM(7443) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7443)))) severity failure;
    assert RAM(7444) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7444)))) severity failure;
    assert RAM(7445) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7445)))) severity failure;
    assert RAM(7446) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7446)))) severity failure;
    assert RAM(7447) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7447)))) severity failure;
    assert RAM(7448) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7448)))) severity failure;
    assert RAM(7449) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7449)))) severity failure;
    assert RAM(7450) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7450)))) severity failure;
    assert RAM(7451) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7451)))) severity failure;
    assert RAM(7452) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7452)))) severity failure;
    assert RAM(7453) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7453)))) severity failure;
    assert RAM(7454) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7454)))) severity failure;
    assert RAM(7455) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7455)))) severity failure;
    assert RAM(7456) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7456)))) severity failure;
    assert RAM(7457) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7457)))) severity failure;
    assert RAM(7458) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7458)))) severity failure;
    assert RAM(7459) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7459)))) severity failure;
    assert RAM(7460) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7460)))) severity failure;
    assert RAM(7461) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7461)))) severity failure;
    assert RAM(7462) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7462)))) severity failure;
    assert RAM(7463) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7463)))) severity failure;
    assert RAM(7464) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7464)))) severity failure;
    assert RAM(7465) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7465)))) severity failure;
    assert RAM(7466) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7466)))) severity failure;
    assert RAM(7467) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7467)))) severity failure;
    assert RAM(7468) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7468)))) severity failure;
    assert RAM(7469) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7469)))) severity failure;
    assert RAM(7470) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7470)))) severity failure;
    assert RAM(7471) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7471)))) severity failure;
    assert RAM(7472) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7472)))) severity failure;
    assert RAM(7473) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7473)))) severity failure;
    assert RAM(7474) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7474)))) severity failure;
    assert RAM(7475) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7475)))) severity failure;
    assert RAM(7476) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7476)))) severity failure;
    assert RAM(7477) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7477)))) severity failure;
    assert RAM(7478) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7478)))) severity failure;
    assert RAM(7479) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7479)))) severity failure;
    assert RAM(7480) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7480)))) severity failure;
    assert RAM(7481) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7481)))) severity failure;
    assert RAM(7482) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7482)))) severity failure;
    assert RAM(7483) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7483)))) severity failure;
    assert RAM(7484) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7484)))) severity failure;
    assert RAM(7485) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7485)))) severity failure;
    assert RAM(7486) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7486)))) severity failure;
    assert RAM(7487) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7487)))) severity failure;
    assert RAM(7488) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7488)))) severity failure;
    assert RAM(7489) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7489)))) severity failure;
    assert RAM(7490) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7490)))) severity failure;
    assert RAM(7491) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7491)))) severity failure;
    assert RAM(7492) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7492)))) severity failure;
    assert RAM(7493) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7493)))) severity failure;
    assert RAM(7494) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7494)))) severity failure;
    assert RAM(7495) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7495)))) severity failure;
    assert RAM(7496) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7496)))) severity failure;
    assert RAM(7497) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7497)))) severity failure;
    assert RAM(7498) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7498)))) severity failure;
    assert RAM(7499) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7499)))) severity failure;
    assert RAM(7500) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7500)))) severity failure;
    assert RAM(7501) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7501)))) severity failure;
    assert RAM(7502) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7502)))) severity failure;
    assert RAM(7503) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7503)))) severity failure;
    assert RAM(7504) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7504)))) severity failure;
    assert RAM(7505) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7505)))) severity failure;
    assert RAM(7506) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7506)))) severity failure;
    assert RAM(7507) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7507)))) severity failure;
    assert RAM(7508) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7508)))) severity failure;
    assert RAM(7509) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7509)))) severity failure;
    assert RAM(7510) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7510)))) severity failure;
    assert RAM(7511) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7511)))) severity failure;
    assert RAM(7512) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7512)))) severity failure;
    assert RAM(7513) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7513)))) severity failure;
    assert RAM(7514) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7514)))) severity failure;
    assert RAM(7515) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7515)))) severity failure;
    assert RAM(7516) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7516)))) severity failure;
    assert RAM(7517) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7517)))) severity failure;
    assert RAM(7518) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7518)))) severity failure;
    assert RAM(7519) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7519)))) severity failure;
    assert RAM(7520) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7520)))) severity failure;
    assert RAM(7521) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7521)))) severity failure;
    assert RAM(7522) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7522)))) severity failure;
    assert RAM(7523) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7523)))) severity failure;
    assert RAM(7524) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7524)))) severity failure;
    assert RAM(7525) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7525)))) severity failure;
    assert RAM(7526) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7526)))) severity failure;
    assert RAM(7527) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7527)))) severity failure;
    assert RAM(7528) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7528)))) severity failure;
    assert RAM(7529) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7529)))) severity failure;
    assert RAM(7530) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7530)))) severity failure;
    assert RAM(7531) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7531)))) severity failure;
    assert RAM(7532) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7532)))) severity failure;
    assert RAM(7533) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7533)))) severity failure;
    assert RAM(7534) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7534)))) severity failure;
    assert RAM(7535) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7535)))) severity failure;
    assert RAM(7536) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7536)))) severity failure;
    assert RAM(7537) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7537)))) severity failure;
    assert RAM(7538) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7538)))) severity failure;
    assert RAM(7539) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7539)))) severity failure;
    assert RAM(7540) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7540)))) severity failure;
    assert RAM(7541) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7541)))) severity failure;
    assert RAM(7542) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7542)))) severity failure;
    assert RAM(7543) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7543)))) severity failure;
    assert RAM(7544) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7544)))) severity failure;
    assert RAM(7545) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7545)))) severity failure;
    assert RAM(7546) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7546)))) severity failure;
    assert RAM(7547) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7547)))) severity failure;
    assert RAM(7548) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7548)))) severity failure;
    assert RAM(7549) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7549)))) severity failure;
    assert RAM(7550) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7550)))) severity failure;
    assert RAM(7551) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7551)))) severity failure;
    assert RAM(7552) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7552)))) severity failure;
    assert RAM(7553) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7553)))) severity failure;
    assert RAM(7554) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7554)))) severity failure;
    assert RAM(7555) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7555)))) severity failure;
    assert RAM(7556) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7556)))) severity failure;
    assert RAM(7557) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7557)))) severity failure;
    assert RAM(7558) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7558)))) severity failure;
    assert RAM(7559) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7559)))) severity failure;
    assert RAM(7560) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7560)))) severity failure;
    assert RAM(7561) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7561)))) severity failure;
    assert RAM(7562) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7562)))) severity failure;
    assert RAM(7563) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7563)))) severity failure;
    assert RAM(7564) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7564)))) severity failure;
    assert RAM(7565) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7565)))) severity failure;
    assert RAM(7566) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7566)))) severity failure;
    assert RAM(7567) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7567)))) severity failure;
    assert RAM(7568) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7568)))) severity failure;
    assert RAM(7569) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7569)))) severity failure;
    assert RAM(7570) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7570)))) severity failure;
    assert RAM(7571) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7571)))) severity failure;
    assert RAM(7572) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7572)))) severity failure;
    assert RAM(7573) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7573)))) severity failure;
    assert RAM(7574) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7574)))) severity failure;
    assert RAM(7575) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7575)))) severity failure;
    assert RAM(7576) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7576)))) severity failure;
    assert RAM(7577) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7577)))) severity failure;
    assert RAM(7578) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7578)))) severity failure;
    assert RAM(7579) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7579)))) severity failure;
    assert RAM(7580) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7580)))) severity failure;
    assert RAM(7581) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7581)))) severity failure;
    assert RAM(7582) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7582)))) severity failure;
    assert RAM(7583) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7583)))) severity failure;
    assert RAM(7584) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7584)))) severity failure;
    assert RAM(7585) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7585)))) severity failure;
    assert RAM(7586) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7586)))) severity failure;
    assert RAM(7587) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7587)))) severity failure;
    assert RAM(7588) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7588)))) severity failure;
    assert RAM(7589) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7589)))) severity failure;
    assert RAM(7590) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7590)))) severity failure;
    assert RAM(7591) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7591)))) severity failure;
    assert RAM(7592) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7592)))) severity failure;
    assert RAM(7593) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7593)))) severity failure;
    assert RAM(7594) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7594)))) severity failure;
    assert RAM(7595) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7595)))) severity failure;
    assert RAM(7596) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7596)))) severity failure;
    assert RAM(7597) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7597)))) severity failure;
    assert RAM(7598) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7598)))) severity failure;
    assert RAM(7599) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7599)))) severity failure;
    assert RAM(7600) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7600)))) severity failure;
    assert RAM(7601) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7601)))) severity failure;
    assert RAM(7602) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7602)))) severity failure;
    assert RAM(7603) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7603)))) severity failure;
    assert RAM(7604) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7604)))) severity failure;
    assert RAM(7605) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7605)))) severity failure;
    assert RAM(7606) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7606)))) severity failure;
    assert RAM(7607) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7607)))) severity failure;
    assert RAM(7608) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7608)))) severity failure;
    assert RAM(7609) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7609)))) severity failure;
    assert RAM(7610) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7610)))) severity failure;
    assert RAM(7611) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7611)))) severity failure;
    assert RAM(7612) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7612)))) severity failure;
    assert RAM(7613) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7613)))) severity failure;
    assert RAM(7614) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7614)))) severity failure;
    assert RAM(7615) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7615)))) severity failure;
    assert RAM(7616) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7616)))) severity failure;
    assert RAM(7617) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7617)))) severity failure;
    assert RAM(7618) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7618)))) severity failure;
    assert RAM(7619) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7619)))) severity failure;
    assert RAM(7620) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7620)))) severity failure;
    assert RAM(7621) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7621)))) severity failure;
    assert RAM(7622) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7622)))) severity failure;
    assert RAM(7623) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7623)))) severity failure;
    assert RAM(7624) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7624)))) severity failure;
    assert RAM(7625) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7625)))) severity failure;
    assert RAM(7626) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7626)))) severity failure;
    assert RAM(7627) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7627)))) severity failure;
    assert RAM(7628) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7628)))) severity failure;
    assert RAM(7629) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7629)))) severity failure;
    assert RAM(7630) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7630)))) severity failure;
    assert RAM(7631) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7631)))) severity failure;
    assert RAM(7632) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7632)))) severity failure;
    assert RAM(7633) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7633)))) severity failure;
    assert RAM(7634) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7634)))) severity failure;
    assert RAM(7635) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7635)))) severity failure;
    assert RAM(7636) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7636)))) severity failure;
    assert RAM(7637) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7637)))) severity failure;
    assert RAM(7638) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7638)))) severity failure;
    assert RAM(7639) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7639)))) severity failure;
    assert RAM(7640) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7640)))) severity failure;
    assert RAM(7641) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7641)))) severity failure;
    assert RAM(7642) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7642)))) severity failure;
    assert RAM(7643) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7643)))) severity failure;
    assert RAM(7644) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7644)))) severity failure;
    assert RAM(7645) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7645)))) severity failure;
    assert RAM(7646) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7646)))) severity failure;
    assert RAM(7647) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7647)))) severity failure;
    assert RAM(7648) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7648)))) severity failure;
    assert RAM(7649) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7649)))) severity failure;
    assert RAM(7650) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7650)))) severity failure;
    assert RAM(7651) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7651)))) severity failure;
    assert RAM(7652) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7652)))) severity failure;
    assert RAM(7653) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7653)))) severity failure;
    assert RAM(7654) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7654)))) severity failure;
    assert RAM(7655) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7655)))) severity failure;
    assert RAM(7656) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7656)))) severity failure;
    assert RAM(7657) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7657)))) severity failure;
    assert RAM(7658) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7658)))) severity failure;
    assert RAM(7659) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7659)))) severity failure;
    assert RAM(7660) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7660)))) severity failure;
    assert RAM(7661) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7661)))) severity failure;
    assert RAM(7662) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7662)))) severity failure;
    assert RAM(7663) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7663)))) severity failure;
    assert RAM(7664) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7664)))) severity failure;
    assert RAM(7665) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7665)))) severity failure;
    assert RAM(7666) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7666)))) severity failure;
    assert RAM(7667) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7667)))) severity failure;
    assert RAM(7668) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7668)))) severity failure;
    assert RAM(7669) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7669)))) severity failure;
    assert RAM(7670) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7670)))) severity failure;
    assert RAM(7671) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7671)))) severity failure;
    assert RAM(7672) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7672)))) severity failure;
    assert RAM(7673) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7673)))) severity failure;
    assert RAM(7674) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7674)))) severity failure;
    assert RAM(7675) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7675)))) severity failure;
    assert RAM(7676) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7676)))) severity failure;
    assert RAM(7677) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7677)))) severity failure;
    assert RAM(7678) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7678)))) severity failure;
    assert RAM(7679) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7679)))) severity failure;
    assert RAM(7680) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7680)))) severity failure;
    assert RAM(7681) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7681)))) severity failure;
    assert RAM(7682) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7682)))) severity failure;
    assert RAM(7683) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7683)))) severity failure;
    assert RAM(7684) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7684)))) severity failure;
    assert RAM(7685) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7685)))) severity failure;
    assert RAM(7686) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7686)))) severity failure;
    assert RAM(7687) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7687)))) severity failure;
    assert RAM(7688) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7688)))) severity failure;
    assert RAM(7689) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7689)))) severity failure;
    assert RAM(7690) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7690)))) severity failure;
    assert RAM(7691) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7691)))) severity failure;
    assert RAM(7692) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7692)))) severity failure;
    assert RAM(7693) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7693)))) severity failure;
    assert RAM(7694) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7694)))) severity failure;
    assert RAM(7695) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7695)))) severity failure;
    assert RAM(7696) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7696)))) severity failure;
    assert RAM(7697) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7697)))) severity failure;
    assert RAM(7698) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7698)))) severity failure;
    assert RAM(7699) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7699)))) severity failure;
    assert RAM(7700) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7700)))) severity failure;
    assert RAM(7701) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7701)))) severity failure;
    assert RAM(7702) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7702)))) severity failure;
    assert RAM(7703) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7703)))) severity failure;
    assert RAM(7704) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7704)))) severity failure;
    assert RAM(7705) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7705)))) severity failure;
    assert RAM(7706) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7706)))) severity failure;
    assert RAM(7707) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7707)))) severity failure;
    assert RAM(7708) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7708)))) severity failure;
    assert RAM(7709) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7709)))) severity failure;
    assert RAM(7710) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7710)))) severity failure;
    assert RAM(7711) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7711)))) severity failure;
    assert RAM(7712) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7712)))) severity failure;
    assert RAM(7713) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7713)))) severity failure;
    assert RAM(7714) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7714)))) severity failure;
    assert RAM(7715) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7715)))) severity failure;
    assert RAM(7716) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7716)))) severity failure;
    assert RAM(7717) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7717)))) severity failure;
    assert RAM(7718) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7718)))) severity failure;
    assert RAM(7719) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7719)))) severity failure;
    assert RAM(7720) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7720)))) severity failure;
    assert RAM(7721) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7721)))) severity failure;
    assert RAM(7722) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7722)))) severity failure;
    assert RAM(7723) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7723)))) severity failure;
    assert RAM(7724) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7724)))) severity failure;
    assert RAM(7725) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7725)))) severity failure;
    assert RAM(7726) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7726)))) severity failure;
    assert RAM(7727) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7727)))) severity failure;
    assert RAM(7728) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7728)))) severity failure;
    assert RAM(7729) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7729)))) severity failure;
    assert RAM(7730) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7730)))) severity failure;
    assert RAM(7731) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7731)))) severity failure;
    assert RAM(7732) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7732)))) severity failure;
    assert RAM(7733) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7733)))) severity failure;
    assert RAM(7734) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7734)))) severity failure;
    assert RAM(7735) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7735)))) severity failure;
    assert RAM(7736) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7736)))) severity failure;
    assert RAM(7737) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7737)))) severity failure;
    assert RAM(7738) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7738)))) severity failure;
    assert RAM(7739) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7739)))) severity failure;
    assert RAM(7740) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7740)))) severity failure;
    assert RAM(7741) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7741)))) severity failure;
    assert RAM(7742) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7742)))) severity failure;
    assert RAM(7743) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7743)))) severity failure;
    assert RAM(7744) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7744)))) severity failure;
    assert RAM(7745) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7745)))) severity failure;
    assert RAM(7746) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7746)))) severity failure;
    assert RAM(7747) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7747)))) severity failure;
    assert RAM(7748) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7748)))) severity failure;
    assert RAM(7749) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7749)))) severity failure;
    assert RAM(7750) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7750)))) severity failure;
    assert RAM(7751) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7751)))) severity failure;
    assert RAM(7752) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7752)))) severity failure;
    assert RAM(7753) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7753)))) severity failure;
    assert RAM(7754) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7754)))) severity failure;
    assert RAM(7755) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7755)))) severity failure;
    assert RAM(7756) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7756)))) severity failure;
    assert RAM(7757) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7757)))) severity failure;
    assert RAM(7758) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7758)))) severity failure;
    assert RAM(7759) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7759)))) severity failure;
    assert RAM(7760) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7760)))) severity failure;
    assert RAM(7761) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7761)))) severity failure;
    assert RAM(7762) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7762)))) severity failure;
    assert RAM(7763) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7763)))) severity failure;
    assert RAM(7764) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7764)))) severity failure;
    assert RAM(7765) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7765)))) severity failure;
    assert RAM(7766) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7766)))) severity failure;
    assert RAM(7767) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7767)))) severity failure;
    assert RAM(7768) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7768)))) severity failure;
    assert RAM(7769) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7769)))) severity failure;
    assert RAM(7770) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7770)))) severity failure;
    assert RAM(7771) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7771)))) severity failure;
    assert RAM(7772) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7772)))) severity failure;
    assert RAM(7773) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7773)))) severity failure;
    assert RAM(7774) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7774)))) severity failure;
    assert RAM(7775) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7775)))) severity failure;
    assert RAM(7776) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7776)))) severity failure;
    assert RAM(7777) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7777)))) severity failure;
    assert RAM(7778) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7778)))) severity failure;
    assert RAM(7779) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7779)))) severity failure;
    assert RAM(7780) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7780)))) severity failure;
    assert RAM(7781) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7781)))) severity failure;
    assert RAM(7782) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7782)))) severity failure;
    assert RAM(7783) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7783)))) severity failure;
    assert RAM(7784) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7784)))) severity failure;
    assert RAM(7785) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7785)))) severity failure;
    assert RAM(7786) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7786)))) severity failure;
    assert RAM(7787) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7787)))) severity failure;
    assert RAM(7788) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7788)))) severity failure;
    assert RAM(7789) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7789)))) severity failure;
    assert RAM(7790) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7790)))) severity failure;
    assert RAM(7791) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7791)))) severity failure;
    assert RAM(7792) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7792)))) severity failure;
    assert RAM(7793) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7793)))) severity failure;
    assert RAM(7794) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7794)))) severity failure;
    assert RAM(7795) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7795)))) severity failure;
    assert RAM(7796) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7796)))) severity failure;
    assert RAM(7797) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7797)))) severity failure;
    assert RAM(7798) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7798)))) severity failure;
    assert RAM(7799) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7799)))) severity failure;
    assert RAM(7800) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7800)))) severity failure;
    assert RAM(7801) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7801)))) severity failure;
    assert RAM(7802) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7802)))) severity failure;
    assert RAM(7803) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7803)))) severity failure;
    assert RAM(7804) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7804)))) severity failure;
    assert RAM(7805) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7805)))) severity failure;
    assert RAM(7806) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7806)))) severity failure;
    assert RAM(7807) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7807)))) severity failure;
    assert RAM(7808) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7808)))) severity failure;
    assert RAM(7809) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7809)))) severity failure;
    assert RAM(7810) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7810)))) severity failure;
    assert RAM(7811) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7811)))) severity failure;
    assert RAM(7812) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7812)))) severity failure;
    assert RAM(7813) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7813)))) severity failure;
    assert RAM(7814) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7814)))) severity failure;
    assert RAM(7815) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7815)))) severity failure;
    assert RAM(7816) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7816)))) severity failure;
    assert RAM(7817) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7817)))) severity failure;
    assert RAM(7818) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7818)))) severity failure;
    assert RAM(7819) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7819)))) severity failure;
    assert RAM(7820) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7820)))) severity failure;
    assert RAM(7821) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7821)))) severity failure;
    assert RAM(7822) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7822)))) severity failure;
    assert RAM(7823) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7823)))) severity failure;
    assert RAM(7824) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7824)))) severity failure;
    assert RAM(7825) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7825)))) severity failure;
    assert RAM(7826) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7826)))) severity failure;
    assert RAM(7827) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7827)))) severity failure;
    assert RAM(7828) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7828)))) severity failure;
    assert RAM(7829) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7829)))) severity failure;
    assert RAM(7830) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7830)))) severity failure;
    assert RAM(7831) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7831)))) severity failure;
    assert RAM(7832) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7832)))) severity failure;
    assert RAM(7833) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7833)))) severity failure;
    assert RAM(7834) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7834)))) severity failure;
    assert RAM(7835) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7835)))) severity failure;
    assert RAM(7836) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7836)))) severity failure;
    assert RAM(7837) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7837)))) severity failure;
    assert RAM(7838) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7838)))) severity failure;
    assert RAM(7839) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7839)))) severity failure;
    assert RAM(7840) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7840)))) severity failure;
    assert RAM(7841) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7841)))) severity failure;
    assert RAM(7842) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7842)))) severity failure;
    assert RAM(7843) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7843)))) severity failure;
    assert RAM(7844) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7844)))) severity failure;
    assert RAM(7845) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7845)))) severity failure;
    assert RAM(7846) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7846)))) severity failure;
    assert RAM(7847) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7847)))) severity failure;
    assert RAM(7848) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7848)))) severity failure;
    assert RAM(7849) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7849)))) severity failure;
    assert RAM(7850) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7850)))) severity failure;
    assert RAM(7851) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7851)))) severity failure;
    assert RAM(7852) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7852)))) severity failure;
    assert RAM(7853) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7853)))) severity failure;
    assert RAM(7854) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7854)))) severity failure;
    assert RAM(7855) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7855)))) severity failure;
    assert RAM(7856) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7856)))) severity failure;
    assert RAM(7857) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7857)))) severity failure;
    assert RAM(7858) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7858)))) severity failure;
    assert RAM(7859) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7859)))) severity failure;
    assert RAM(7860) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7860)))) severity failure;
    assert RAM(7861) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7861)))) severity failure;
    assert RAM(7862) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7862)))) severity failure;
    assert RAM(7863) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7863)))) severity failure;
    assert RAM(7864) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7864)))) severity failure;
    assert RAM(7865) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7865)))) severity failure;
    assert RAM(7866) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7866)))) severity failure;
    assert RAM(7867) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7867)))) severity failure;
    assert RAM(7868) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7868)))) severity failure;
    assert RAM(7869) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7869)))) severity failure;
    assert RAM(7870) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7870)))) severity failure;
    assert RAM(7871) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7871)))) severity failure;
    assert RAM(7872) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7872)))) severity failure;
    assert RAM(7873) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7873)))) severity failure;
    assert RAM(7874) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7874)))) severity failure;
    assert RAM(7875) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7875)))) severity failure;
    assert RAM(7876) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7876)))) severity failure;
    assert RAM(7877) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7877)))) severity failure;
    assert RAM(7878) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7878)))) severity failure;
    assert RAM(7879) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7879)))) severity failure;
    assert RAM(7880) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7880)))) severity failure;
    assert RAM(7881) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7881)))) severity failure;
    assert RAM(7882) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7882)))) severity failure;
    assert RAM(7883) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7883)))) severity failure;
    assert RAM(7884) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7884)))) severity failure;
    assert RAM(7885) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7885)))) severity failure;
    assert RAM(7886) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7886)))) severity failure;
    assert RAM(7887) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7887)))) severity failure;
    assert RAM(7888) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7888)))) severity failure;
    assert RAM(7889) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7889)))) severity failure;
    assert RAM(7890) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7890)))) severity failure;
    assert RAM(7891) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7891)))) severity failure;
    assert RAM(7892) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7892)))) severity failure;
    assert RAM(7893) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7893)))) severity failure;
    assert RAM(7894) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7894)))) severity failure;
    assert RAM(7895) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7895)))) severity failure;
    assert RAM(7896) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7896)))) severity failure;
    assert RAM(7897) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7897)))) severity failure;
    assert RAM(7898) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7898)))) severity failure;
    assert RAM(7899) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7899)))) severity failure;
    assert RAM(7900) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7900)))) severity failure;
    assert RAM(7901) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7901)))) severity failure;
    assert RAM(7902) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7902)))) severity failure;
    assert RAM(7903) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7903)))) severity failure;
    assert RAM(7904) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7904)))) severity failure;
    assert RAM(7905) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7905)))) severity failure;
    assert RAM(7906) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7906)))) severity failure;
    assert RAM(7907) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7907)))) severity failure;
    assert RAM(7908) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7908)))) severity failure;
    assert RAM(7909) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7909)))) severity failure;
    assert RAM(7910) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7910)))) severity failure;
    assert RAM(7911) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7911)))) severity failure;
    assert RAM(7912) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7912)))) severity failure;
    assert RAM(7913) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7913)))) severity failure;
    assert RAM(7914) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7914)))) severity failure;
    assert RAM(7915) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7915)))) severity failure;
    assert RAM(7916) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7916)))) severity failure;
    assert RAM(7917) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7917)))) severity failure;
    assert RAM(7918) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7918)))) severity failure;
    assert RAM(7919) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7919)))) severity failure;
    assert RAM(7920) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7920)))) severity failure;
    assert RAM(7921) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7921)))) severity failure;
    assert RAM(7922) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7922)))) severity failure;
    assert RAM(7923) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7923)))) severity failure;
    assert RAM(7924) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7924)))) severity failure;
    assert RAM(7925) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7925)))) severity failure;
    assert RAM(7926) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7926)))) severity failure;
    assert RAM(7927) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7927)))) severity failure;
    assert RAM(7928) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7928)))) severity failure;
    assert RAM(7929) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7929)))) severity failure;
    assert RAM(7930) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7930)))) severity failure;
    assert RAM(7931) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7931)))) severity failure;
    assert RAM(7932) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7932)))) severity failure;
    assert RAM(7933) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7933)))) severity failure;
    assert RAM(7934) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7934)))) severity failure;
    assert RAM(7935) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7935)))) severity failure;
    assert RAM(7936) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7936)))) severity failure;
    assert RAM(7937) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7937)))) severity failure;
    assert RAM(7938) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7938)))) severity failure;
    assert RAM(7939) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7939)))) severity failure;
    assert RAM(7940) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7940)))) severity failure;
    assert RAM(7941) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7941)))) severity failure;
    assert RAM(7942) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7942)))) severity failure;
    assert RAM(7943) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7943)))) severity failure;
    assert RAM(7944) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7944)))) severity failure;
    assert RAM(7945) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7945)))) severity failure;
    assert RAM(7946) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7946)))) severity failure;
    assert RAM(7947) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7947)))) severity failure;
    assert RAM(7948) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7948)))) severity failure;
    assert RAM(7949) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7949)))) severity failure;
    assert RAM(7950) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7950)))) severity failure;
    assert RAM(7951) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7951)))) severity failure;
    assert RAM(7952) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7952)))) severity failure;
    assert RAM(7953) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7953)))) severity failure;
    assert RAM(7954) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7954)))) severity failure;
    assert RAM(7955) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7955)))) severity failure;
    assert RAM(7956) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7956)))) severity failure;
    assert RAM(7957) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7957)))) severity failure;
    assert RAM(7958) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7958)))) severity failure;
    assert RAM(7959) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7959)))) severity failure;
    assert RAM(7960) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7960)))) severity failure;
    assert RAM(7961) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7961)))) severity failure;
    assert RAM(7962) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7962)))) severity failure;
    assert RAM(7963) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7963)))) severity failure;
    assert RAM(7964) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7964)))) severity failure;
    assert RAM(7965) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7965)))) severity failure;
    assert RAM(7966) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7966)))) severity failure;
    assert RAM(7967) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7967)))) severity failure;
    assert RAM(7968) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7968)))) severity failure;
    assert RAM(7969) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7969)))) severity failure;
    assert RAM(7970) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7970)))) severity failure;
    assert RAM(7971) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7971)))) severity failure;
    assert RAM(7972) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7972)))) severity failure;
    assert RAM(7973) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7973)))) severity failure;
    assert RAM(7974) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7974)))) severity failure;
    assert RAM(7975) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7975)))) severity failure;
    assert RAM(7976) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7976)))) severity failure;
    assert RAM(7977) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7977)))) severity failure;
    assert RAM(7978) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7978)))) severity failure;
    assert RAM(7979) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7979)))) severity failure;
    assert RAM(7980) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7980)))) severity failure;
    assert RAM(7981) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7981)))) severity failure;
    assert RAM(7982) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7982)))) severity failure;
    assert RAM(7983) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7983)))) severity failure;
    assert RAM(7984) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7984)))) severity failure;
    assert RAM(7985) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7985)))) severity failure;
    assert RAM(7986) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7986)))) severity failure;
    assert RAM(7987) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7987)))) severity failure;
    assert RAM(7988) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7988)))) severity failure;
    assert RAM(7989) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7989)))) severity failure;
    assert RAM(7990) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7990)))) severity failure;
    assert RAM(7991) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7991)))) severity failure;
    assert RAM(7992) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7992)))) severity failure;
    assert RAM(7993) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7993)))) severity failure;
    assert RAM(7994) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7994)))) severity failure;
    assert RAM(7995) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7995)))) severity failure;
    assert RAM(7996) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7996)))) severity failure;
    assert RAM(7997) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7997)))) severity failure;
    assert RAM(7998) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(7998)))) severity failure;
    assert RAM(7999) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(7999)))) severity failure;
    assert RAM(8000) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8000)))) severity failure;
    assert RAM(8001) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8001)))) severity failure;
    assert RAM(8002) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8002)))) severity failure;
    assert RAM(8003) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8003)))) severity failure;
    assert RAM(8004) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8004)))) severity failure;
    assert RAM(8005) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8005)))) severity failure;
    assert RAM(8006) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8006)))) severity failure;
    assert RAM(8007) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8007)))) severity failure;
    assert RAM(8008) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8008)))) severity failure;
    assert RAM(8009) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8009)))) severity failure;
    assert RAM(8010) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8010)))) severity failure;
    assert RAM(8011) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8011)))) severity failure;
    assert RAM(8012) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8012)))) severity failure;
    assert RAM(8013) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8013)))) severity failure;
    assert RAM(8014) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8014)))) severity failure;
    assert RAM(8015) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8015)))) severity failure;
    assert RAM(8016) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8016)))) severity failure;
    assert RAM(8017) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8017)))) severity failure;
    assert RAM(8018) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8018)))) severity failure;
    assert RAM(8019) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8019)))) severity failure;
    assert RAM(8020) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8020)))) severity failure;
    assert RAM(8021) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8021)))) severity failure;
    assert RAM(8022) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8022)))) severity failure;
    assert RAM(8023) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8023)))) severity failure;
    assert RAM(8024) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8024)))) severity failure;
    assert RAM(8025) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8025)))) severity failure;
    assert RAM(8026) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8026)))) severity failure;
    assert RAM(8027) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8027)))) severity failure;
    assert RAM(8028) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8028)))) severity failure;
    assert RAM(8029) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8029)))) severity failure;
    assert RAM(8030) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8030)))) severity failure;
    assert RAM(8031) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8031)))) severity failure;
    assert RAM(8032) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8032)))) severity failure;
    assert RAM(8033) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8033)))) severity failure;
    assert RAM(8034) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8034)))) severity failure;
    assert RAM(8035) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8035)))) severity failure;
    assert RAM(8036) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8036)))) severity failure;
    assert RAM(8037) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8037)))) severity failure;
    assert RAM(8038) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8038)))) severity failure;
    assert RAM(8039) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8039)))) severity failure;
    assert RAM(8040) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8040)))) severity failure;
    assert RAM(8041) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8041)))) severity failure;
    assert RAM(8042) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8042)))) severity failure;
    assert RAM(8043) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8043)))) severity failure;
    assert RAM(8044) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8044)))) severity failure;
    assert RAM(8045) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8045)))) severity failure;
    assert RAM(8046) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8046)))) severity failure;
    assert RAM(8047) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8047)))) severity failure;
    assert RAM(8048) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8048)))) severity failure;
    assert RAM(8049) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8049)))) severity failure;
    assert RAM(8050) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8050)))) severity failure;
    assert RAM(8051) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8051)))) severity failure;
    assert RAM(8052) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8052)))) severity failure;
    assert RAM(8053) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8053)))) severity failure;
    assert RAM(8054) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8054)))) severity failure;
    assert RAM(8055) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8055)))) severity failure;
    assert RAM(8056) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8056)))) severity failure;
    assert RAM(8057) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8057)))) severity failure;
    assert RAM(8058) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8058)))) severity failure;
    assert RAM(8059) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8059)))) severity failure;
    assert RAM(8060) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8060)))) severity failure;
    assert RAM(8061) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8061)))) severity failure;
    assert RAM(8062) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8062)))) severity failure;
    assert RAM(8063) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8063)))) severity failure;
    assert RAM(8064) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8064)))) severity failure;
    assert RAM(8065) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8065)))) severity failure;
    assert RAM(8066) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8066)))) severity failure;
    assert RAM(8067) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8067)))) severity failure;
    assert RAM(8068) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8068)))) severity failure;
    assert RAM(8069) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8069)))) severity failure;
    assert RAM(8070) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8070)))) severity failure;
    assert RAM(8071) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8071)))) severity failure;
    assert RAM(8072) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8072)))) severity failure;
    assert RAM(8073) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8073)))) severity failure;
    assert RAM(8074) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8074)))) severity failure;
    assert RAM(8075) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8075)))) severity failure;
    assert RAM(8076) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8076)))) severity failure;
    assert RAM(8077) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8077)))) severity failure;
    assert RAM(8078) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8078)))) severity failure;
    assert RAM(8079) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8079)))) severity failure;
    assert RAM(8080) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8080)))) severity failure;
    assert RAM(8081) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8081)))) severity failure;
    assert RAM(8082) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8082)))) severity failure;
    assert RAM(8083) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8083)))) severity failure;
    assert RAM(8084) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8084)))) severity failure;
    assert RAM(8085) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8085)))) severity failure;
    assert RAM(8086) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8086)))) severity failure;
    assert RAM(8087) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8087)))) severity failure;
    assert RAM(8088) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8088)))) severity failure;
    assert RAM(8089) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8089)))) severity failure;
    assert RAM(8090) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8090)))) severity failure;
    assert RAM(8091) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8091)))) severity failure;
    assert RAM(8092) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8092)))) severity failure;
    assert RAM(8093) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8093)))) severity failure;
    assert RAM(8094) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8094)))) severity failure;
    assert RAM(8095) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8095)))) severity failure;
    assert RAM(8096) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8096)))) severity failure;
    assert RAM(8097) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8097)))) severity failure;
    assert RAM(8098) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8098)))) severity failure;
    assert RAM(8099) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8099)))) severity failure;
    assert RAM(8100) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8100)))) severity failure;
    assert RAM(8101) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8101)))) severity failure;
    assert RAM(8102) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8102)))) severity failure;
    assert RAM(8103) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8103)))) severity failure;
    assert RAM(8104) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8104)))) severity failure;
    assert RAM(8105) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8105)))) severity failure;
    assert RAM(8106) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8106)))) severity failure;
    assert RAM(8107) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8107)))) severity failure;
    assert RAM(8108) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8108)))) severity failure;
    assert RAM(8109) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8109)))) severity failure;
    assert RAM(8110) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8110)))) severity failure;
    assert RAM(8111) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8111)))) severity failure;
    assert RAM(8112) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8112)))) severity failure;
    assert RAM(8113) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8113)))) severity failure;
    assert RAM(8114) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8114)))) severity failure;
    assert RAM(8115) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8115)))) severity failure;
    assert RAM(8116) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8116)))) severity failure;
    assert RAM(8117) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8117)))) severity failure;
    assert RAM(8118) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8118)))) severity failure;
    assert RAM(8119) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8119)))) severity failure;
    assert RAM(8120) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8120)))) severity failure;
    assert RAM(8121) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8121)))) severity failure;
    assert RAM(8122) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8122)))) severity failure;
    assert RAM(8123) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8123)))) severity failure;
    assert RAM(8124) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8124)))) severity failure;
    assert RAM(8125) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8125)))) severity failure;
    assert RAM(8126) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8126)))) severity failure;
    assert RAM(8127) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8127)))) severity failure;
    assert RAM(8128) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8128)))) severity failure;
    assert RAM(8129) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8129)))) severity failure;
    assert RAM(8130) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8130)))) severity failure;
    assert RAM(8131) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8131)))) severity failure;
    assert RAM(8132) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8132)))) severity failure;
    assert RAM(8133) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8133)))) severity failure;
    assert RAM(8134) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8134)))) severity failure;
    assert RAM(8135) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8135)))) severity failure;
    assert RAM(8136) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8136)))) severity failure;
    assert RAM(8137) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8137)))) severity failure;
    assert RAM(8138) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8138)))) severity failure;
    assert RAM(8139) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8139)))) severity failure;
    assert RAM(8140) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8140)))) severity failure;
    assert RAM(8141) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8141)))) severity failure;
    assert RAM(8142) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8142)))) severity failure;
    assert RAM(8143) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8143)))) severity failure;
    assert RAM(8144) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8144)))) severity failure;
    assert RAM(8145) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8145)))) severity failure;
    assert RAM(8146) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8146)))) severity failure;
    assert RAM(8147) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8147)))) severity failure;
    assert RAM(8148) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8148)))) severity failure;
    assert RAM(8149) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8149)))) severity failure;
    assert RAM(8150) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8150)))) severity failure;
    assert RAM(8151) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8151)))) severity failure;
    assert RAM(8152) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8152)))) severity failure;
    assert RAM(8153) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8153)))) severity failure;
    assert RAM(8154) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8154)))) severity failure;
    assert RAM(8155) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8155)))) severity failure;
    assert RAM(8156) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8156)))) severity failure;
    assert RAM(8157) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8157)))) severity failure;
    assert RAM(8158) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8158)))) severity failure;
    assert RAM(8159) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8159)))) severity failure;
    assert RAM(8160) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8160)))) severity failure;
    assert RAM(8161) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8161)))) severity failure;
    assert RAM(8162) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8162)))) severity failure;
    assert RAM(8163) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8163)))) severity failure;
    assert RAM(8164) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8164)))) severity failure;
    assert RAM(8165) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8165)))) severity failure;
    assert RAM(8166) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8166)))) severity failure;
    assert RAM(8167) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8167)))) severity failure;
    assert RAM(8168) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8168)))) severity failure;
    assert RAM(8169) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8169)))) severity failure;
    assert RAM(8170) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8170)))) severity failure;
    assert RAM(8171) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8171)))) severity failure;
    assert RAM(8172) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8172)))) severity failure;
    assert RAM(8173) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8173)))) severity failure;
    assert RAM(8174) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8174)))) severity failure;
    assert RAM(8175) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8175)))) severity failure;
    assert RAM(8176) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8176)))) severity failure;
    assert RAM(8177) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8177)))) severity failure;
    assert RAM(8178) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8178)))) severity failure;
    assert RAM(8179) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8179)))) severity failure;
    assert RAM(8180) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8180)))) severity failure;
    assert RAM(8181) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8181)))) severity failure;
    assert RAM(8182) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8182)))) severity failure;
    assert RAM(8183) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8183)))) severity failure;
    assert RAM(8184) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8184)))) severity failure;
    assert RAM(8185) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8185)))) severity failure;
    assert RAM(8186) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8186)))) severity failure;
    assert RAM(8187) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8187)))) severity failure;
    assert RAM(8188) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8188)))) severity failure;
    assert RAM(8189) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8189)))) severity failure;
    assert RAM(8190) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8190)))) severity failure;
    assert RAM(8191) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8191)))) severity failure;
    assert RAM(8192) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8192)))) severity failure;
    assert RAM(8193) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8193)))) severity failure;
    assert RAM(8194) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8194)))) severity failure;
    assert RAM(8195) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8195)))) severity failure;
    assert RAM(8196) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8196)))) severity failure;
    assert RAM(8197) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8197)))) severity failure;
    assert RAM(8198) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8198)))) severity failure;
    assert RAM(8199) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8199)))) severity failure;
    assert RAM(8200) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8200)))) severity failure;
    assert RAM(8201) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8201)))) severity failure;
    assert RAM(8202) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8202)))) severity failure;
    assert RAM(8203) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8203)))) severity failure;
    assert RAM(8204) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8204)))) severity failure;
    assert RAM(8205) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8205)))) severity failure;
    assert RAM(8206) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8206)))) severity failure;
    assert RAM(8207) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8207)))) severity failure;
    assert RAM(8208) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8208)))) severity failure;
    assert RAM(8209) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8209)))) severity failure;
    assert RAM(8210) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8210)))) severity failure;
    assert RAM(8211) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8211)))) severity failure;
    assert RAM(8212) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8212)))) severity failure;
    assert RAM(8213) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8213)))) severity failure;
    assert RAM(8214) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8214)))) severity failure;
    assert RAM(8215) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8215)))) severity failure;
    assert RAM(8216) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8216)))) severity failure;
    assert RAM(8217) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8217)))) severity failure;
    assert RAM(8218) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8218)))) severity failure;
    assert RAM(8219) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8219)))) severity failure;
    assert RAM(8220) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8220)))) severity failure;
    assert RAM(8221) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8221)))) severity failure;
    assert RAM(8222) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8222)))) severity failure;
    assert RAM(8223) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8223)))) severity failure;
    assert RAM(8224) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8224)))) severity failure;
    assert RAM(8225) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8225)))) severity failure;
    assert RAM(8226) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8226)))) severity failure;
    assert RAM(8227) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8227)))) severity failure;
    assert RAM(8228) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8228)))) severity failure;
    assert RAM(8229) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8229)))) severity failure;
    assert RAM(8230) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8230)))) severity failure;
    assert RAM(8231) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8231)))) severity failure;
    assert RAM(8232) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8232)))) severity failure;
    assert RAM(8233) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8233)))) severity failure;
    assert RAM(8234) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8234)))) severity failure;
    assert RAM(8235) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8235)))) severity failure;
    assert RAM(8236) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8236)))) severity failure;
    assert RAM(8237) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8237)))) severity failure;
    assert RAM(8238) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8238)))) severity failure;
    assert RAM(8239) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8239)))) severity failure;
    assert RAM(8240) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8240)))) severity failure;
    assert RAM(8241) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8241)))) severity failure;
    assert RAM(8242) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8242)))) severity failure;
    assert RAM(8243) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8243)))) severity failure;
    assert RAM(8244) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8244)))) severity failure;
    assert RAM(8245) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8245)))) severity failure;
    assert RAM(8246) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8246)))) severity failure;
    assert RAM(8247) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8247)))) severity failure;
    assert RAM(8248) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8248)))) severity failure;
    assert RAM(8249) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8249)))) severity failure;
    assert RAM(8250) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8250)))) severity failure;
    assert RAM(8251) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8251)))) severity failure;
    assert RAM(8252) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8252)))) severity failure;
    assert RAM(8253) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8253)))) severity failure;
    assert RAM(8254) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8254)))) severity failure;
    assert RAM(8255) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8255)))) severity failure;
    assert RAM(8256) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8256)))) severity failure;
    assert RAM(8257) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8257)))) severity failure;
    assert RAM(8258) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8258)))) severity failure;
    assert RAM(8259) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8259)))) severity failure;
    assert RAM(8260) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8260)))) severity failure;
    assert RAM(8261) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8261)))) severity failure;
    assert RAM(8262) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8262)))) severity failure;
    assert RAM(8263) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8263)))) severity failure;
    assert RAM(8264) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8264)))) severity failure;
    assert RAM(8265) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8265)))) severity failure;
    assert RAM(8266) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8266)))) severity failure;
    assert RAM(8267) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8267)))) severity failure;
    assert RAM(8268) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8268)))) severity failure;
    assert RAM(8269) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8269)))) severity failure;
    assert RAM(8270) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8270)))) severity failure;
    assert RAM(8271) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8271)))) severity failure;
    assert RAM(8272) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8272)))) severity failure;
    assert RAM(8273) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8273)))) severity failure;
    assert RAM(8274) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8274)))) severity failure;
    assert RAM(8275) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8275)))) severity failure;
    assert RAM(8276) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8276)))) severity failure;
    assert RAM(8277) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8277)))) severity failure;
    assert RAM(8278) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8278)))) severity failure;
    assert RAM(8279) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8279)))) severity failure;
    assert RAM(8280) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8280)))) severity failure;
    assert RAM(8281) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8281)))) severity failure;
    assert RAM(8282) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8282)))) severity failure;
    assert RAM(8283) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8283)))) severity failure;
    assert RAM(8284) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8284)))) severity failure;
    assert RAM(8285) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8285)))) severity failure;
    assert RAM(8286) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8286)))) severity failure;
    assert RAM(8287) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8287)))) severity failure;
    assert RAM(8288) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8288)))) severity failure;
    assert RAM(8289) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8289)))) severity failure;
    assert RAM(8290) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8290)))) severity failure;
    assert RAM(8291) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8291)))) severity failure;
    assert RAM(8292) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8292)))) severity failure;
    assert RAM(8293) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8293)))) severity failure;
    assert RAM(8294) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8294)))) severity failure;
    assert RAM(8295) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8295)))) severity failure;
    assert RAM(8296) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8296)))) severity failure;
    assert RAM(8297) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8297)))) severity failure;
    assert RAM(8298) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8298)))) severity failure;
    assert RAM(8299) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8299)))) severity failure;
    assert RAM(8300) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8300)))) severity failure;
    assert RAM(8301) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8301)))) severity failure;
    assert RAM(8302) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8302)))) severity failure;
    assert RAM(8303) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8303)))) severity failure;
    assert RAM(8304) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8304)))) severity failure;
    assert RAM(8305) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8305)))) severity failure;
    assert RAM(8306) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8306)))) severity failure;
    assert RAM(8307) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8307)))) severity failure;
    assert RAM(8308) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8308)))) severity failure;
    assert RAM(8309) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8309)))) severity failure;
    assert RAM(8310) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8310)))) severity failure;
    assert RAM(8311) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8311)))) severity failure;
    assert RAM(8312) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8312)))) severity failure;
    assert RAM(8313) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8313)))) severity failure;
    assert RAM(8314) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8314)))) severity failure;
    assert RAM(8315) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8315)))) severity failure;
    assert RAM(8316) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8316)))) severity failure;
    assert RAM(8317) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8317)))) severity failure;
    assert RAM(8318) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8318)))) severity failure;
    assert RAM(8319) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8319)))) severity failure;
    assert RAM(8320) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8320)))) severity failure;
    assert RAM(8321) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8321)))) severity failure;
    assert RAM(8322) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8322)))) severity failure;
    assert RAM(8323) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8323)))) severity failure;
    assert RAM(8324) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8324)))) severity failure;
    assert RAM(8325) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8325)))) severity failure;
    assert RAM(8326) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8326)))) severity failure;
    assert RAM(8327) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8327)))) severity failure;
    assert RAM(8328) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8328)))) severity failure;
    assert RAM(8329) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8329)))) severity failure;
    assert RAM(8330) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8330)))) severity failure;
    assert RAM(8331) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8331)))) severity failure;
    assert RAM(8332) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8332)))) severity failure;
    assert RAM(8333) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8333)))) severity failure;
    assert RAM(8334) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8334)))) severity failure;
    assert RAM(8335) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8335)))) severity failure;
    assert RAM(8336) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8336)))) severity failure;
    assert RAM(8337) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8337)))) severity failure;
    assert RAM(8338) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8338)))) severity failure;
    assert RAM(8339) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8339)))) severity failure;
    assert RAM(8340) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8340)))) severity failure;
    assert RAM(8341) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8341)))) severity failure;
    assert RAM(8342) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8342)))) severity failure;
    assert RAM(8343) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8343)))) severity failure;
    assert RAM(8344) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8344)))) severity failure;
    assert RAM(8345) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8345)))) severity failure;
    assert RAM(8346) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8346)))) severity failure;
    assert RAM(8347) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8347)))) severity failure;
    assert RAM(8348) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8348)))) severity failure;
    assert RAM(8349) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8349)))) severity failure;
    assert RAM(8350) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8350)))) severity failure;
    assert RAM(8351) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8351)))) severity failure;
    assert RAM(8352) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8352)))) severity failure;
    assert RAM(8353) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8353)))) severity failure;
    assert RAM(8354) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8354)))) severity failure;
    assert RAM(8355) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8355)))) severity failure;
    assert RAM(8356) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8356)))) severity failure;
    assert RAM(8357) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8357)))) severity failure;
    assert RAM(8358) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8358)))) severity failure;
    assert RAM(8359) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8359)))) severity failure;
    assert RAM(8360) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8360)))) severity failure;
    assert RAM(8361) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8361)))) severity failure;
    assert RAM(8362) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8362)))) severity failure;
    assert RAM(8363) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8363)))) severity failure;
    assert RAM(8364) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8364)))) severity failure;
    assert RAM(8365) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8365)))) severity failure;
    assert RAM(8366) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8366)))) severity failure;
    assert RAM(8367) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8367)))) severity failure;
    assert RAM(8368) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8368)))) severity failure;
    assert RAM(8369) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8369)))) severity failure;
    assert RAM(8370) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8370)))) severity failure;
    assert RAM(8371) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8371)))) severity failure;
    assert RAM(8372) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8372)))) severity failure;
    assert RAM(8373) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8373)))) severity failure;
    assert RAM(8374) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8374)))) severity failure;
    assert RAM(8375) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8375)))) severity failure;
    assert RAM(8376) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8376)))) severity failure;
    assert RAM(8377) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8377)))) severity failure;
    assert RAM(8378) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8378)))) severity failure;
    assert RAM(8379) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8379)))) severity failure;
    assert RAM(8380) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8380)))) severity failure;
    assert RAM(8381) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8381)))) severity failure;
    assert RAM(8382) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8382)))) severity failure;
    assert RAM(8383) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8383)))) severity failure;
    assert RAM(8384) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8384)))) severity failure;
    assert RAM(8385) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8385)))) severity failure;
    assert RAM(8386) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8386)))) severity failure;
    assert RAM(8387) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8387)))) severity failure;
    assert RAM(8388) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8388)))) severity failure;
    assert RAM(8389) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8389)))) severity failure;
    assert RAM(8390) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8390)))) severity failure;
    assert RAM(8391) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8391)))) severity failure;
    assert RAM(8392) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8392)))) severity failure;
    assert RAM(8393) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8393)))) severity failure;
    assert RAM(8394) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8394)))) severity failure;
    assert RAM(8395) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8395)))) severity failure;
    assert RAM(8396) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8396)))) severity failure;
    assert RAM(8397) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8397)))) severity failure;
    assert RAM(8398) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8398)))) severity failure;
    assert RAM(8399) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8399)))) severity failure;
    assert RAM(8400) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8400)))) severity failure;
    assert RAM(8401) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8401)))) severity failure;
    assert RAM(8402) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8402)))) severity failure;
    assert RAM(8403) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8403)))) severity failure;
    assert RAM(8404) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8404)))) severity failure;
    assert RAM(8405) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8405)))) severity failure;
    assert RAM(8406) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8406)))) severity failure;
    assert RAM(8407) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8407)))) severity failure;
    assert RAM(8408) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8408)))) severity failure;
    assert RAM(8409) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8409)))) severity failure;
    assert RAM(8410) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8410)))) severity failure;
    assert RAM(8411) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8411)))) severity failure;
    assert RAM(8412) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8412)))) severity failure;
    assert RAM(8413) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8413)))) severity failure;
    assert RAM(8414) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8414)))) severity failure;
    assert RAM(8415) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8415)))) severity failure;
    assert RAM(8416) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8416)))) severity failure;
    assert RAM(8417) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8417)))) severity failure;
    assert RAM(8418) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8418)))) severity failure;
    assert RAM(8419) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8419)))) severity failure;
    assert RAM(8420) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8420)))) severity failure;
    assert RAM(8421) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8421)))) severity failure;
    assert RAM(8422) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8422)))) severity failure;
    assert RAM(8423) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8423)))) severity failure;
    assert RAM(8424) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8424)))) severity failure;
    assert RAM(8425) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8425)))) severity failure;
    assert RAM(8426) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8426)))) severity failure;
    assert RAM(8427) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8427)))) severity failure;
    assert RAM(8428) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8428)))) severity failure;
    assert RAM(8429) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8429)))) severity failure;
    assert RAM(8430) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8430)))) severity failure;
    assert RAM(8431) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8431)))) severity failure;
    assert RAM(8432) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8432)))) severity failure;
    assert RAM(8433) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8433)))) severity failure;
    assert RAM(8434) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8434)))) severity failure;
    assert RAM(8435) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8435)))) severity failure;
    assert RAM(8436) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8436)))) severity failure;
    assert RAM(8437) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8437)))) severity failure;
    assert RAM(8438) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8438)))) severity failure;
    assert RAM(8439) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8439)))) severity failure;
    assert RAM(8440) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8440)))) severity failure;
    assert RAM(8441) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8441)))) severity failure;
    assert RAM(8442) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8442)))) severity failure;
    assert RAM(8443) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8443)))) severity failure;
    assert RAM(8444) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8444)))) severity failure;
    assert RAM(8445) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8445)))) severity failure;
    assert RAM(8446) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8446)))) severity failure;
    assert RAM(8447) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8447)))) severity failure;
    assert RAM(8448) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8448)))) severity failure;
    assert RAM(8449) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8449)))) severity failure;
    assert RAM(8450) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8450)))) severity failure;
    assert RAM(8451) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8451)))) severity failure;
    assert RAM(8452) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8452)))) severity failure;
    assert RAM(8453) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8453)))) severity failure;
    assert RAM(8454) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8454)))) severity failure;
    assert RAM(8455) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8455)))) severity failure;
    assert RAM(8456) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8456)))) severity failure;
    assert RAM(8457) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8457)))) severity failure;
    assert RAM(8458) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8458)))) severity failure;
    assert RAM(8459) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8459)))) severity failure;
    assert RAM(8460) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8460)))) severity failure;
    assert RAM(8461) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8461)))) severity failure;
    assert RAM(8462) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8462)))) severity failure;
    assert RAM(8463) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8463)))) severity failure;
    assert RAM(8464) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8464)))) severity failure;
    assert RAM(8465) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8465)))) severity failure;
    assert RAM(8466) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8466)))) severity failure;
    assert RAM(8467) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8467)))) severity failure;
    assert RAM(8468) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8468)))) severity failure;
    assert RAM(8469) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8469)))) severity failure;
    assert RAM(8470) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8470)))) severity failure;
    assert RAM(8471) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8471)))) severity failure;
    assert RAM(8472) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8472)))) severity failure;
    assert RAM(8473) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8473)))) severity failure;
    assert RAM(8474) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8474)))) severity failure;
    assert RAM(8475) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8475)))) severity failure;
    assert RAM(8476) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8476)))) severity failure;
    assert RAM(8477) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8477)))) severity failure;
    assert RAM(8478) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8478)))) severity failure;
    assert RAM(8479) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8479)))) severity failure;
    assert RAM(8480) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8480)))) severity failure;
    assert RAM(8481) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8481)))) severity failure;
    assert RAM(8482) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8482)))) severity failure;
    assert RAM(8483) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8483)))) severity failure;
    assert RAM(8484) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8484)))) severity failure;
    assert RAM(8485) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8485)))) severity failure;
    assert RAM(8486) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8486)))) severity failure;
    assert RAM(8487) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8487)))) severity failure;
    assert RAM(8488) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8488)))) severity failure;
    assert RAM(8489) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8489)))) severity failure;
    assert RAM(8490) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8490)))) severity failure;
    assert RAM(8491) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8491)))) severity failure;
    assert RAM(8492) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8492)))) severity failure;
    assert RAM(8493) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8493)))) severity failure;
    assert RAM(8494) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8494)))) severity failure;
    assert RAM(8495) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8495)))) severity failure;
    assert RAM(8496) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8496)))) severity failure;
    assert RAM(8497) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8497)))) severity failure;
    assert RAM(8498) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8498)))) severity failure;
    assert RAM(8499) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8499)))) severity failure;
    assert RAM(8500) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8500)))) severity failure;
    assert RAM(8501) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8501)))) severity failure;
    assert RAM(8502) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8502)))) severity failure;
    assert RAM(8503) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8503)))) severity failure;
    assert RAM(8504) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8504)))) severity failure;
    assert RAM(8505) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8505)))) severity failure;
    assert RAM(8506) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8506)))) severity failure;
    assert RAM(8507) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8507)))) severity failure;
    assert RAM(8508) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8508)))) severity failure;
    assert RAM(8509) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8509)))) severity failure;
    assert RAM(8510) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8510)))) severity failure;
    assert RAM(8511) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8511)))) severity failure;
    assert RAM(8512) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8512)))) severity failure;
    assert RAM(8513) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8513)))) severity failure;
    assert RAM(8514) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8514)))) severity failure;
    assert RAM(8515) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8515)))) severity failure;
    assert RAM(8516) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8516)))) severity failure;
    assert RAM(8517) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8517)))) severity failure;
    assert RAM(8518) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8518)))) severity failure;
    assert RAM(8519) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8519)))) severity failure;
    assert RAM(8520) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8520)))) severity failure;
    assert RAM(8521) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8521)))) severity failure;
    assert RAM(8522) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8522)))) severity failure;
    assert RAM(8523) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8523)))) severity failure;
    assert RAM(8524) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8524)))) severity failure;
    assert RAM(8525) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8525)))) severity failure;
    assert RAM(8526) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8526)))) severity failure;
    assert RAM(8527) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8527)))) severity failure;
    assert RAM(8528) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8528)))) severity failure;
    assert RAM(8529) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8529)))) severity failure;
    assert RAM(8530) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8530)))) severity failure;
    assert RAM(8531) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8531)))) severity failure;
    assert RAM(8532) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8532)))) severity failure;
    assert RAM(8533) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8533)))) severity failure;
    assert RAM(8534) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8534)))) severity failure;
    assert RAM(8535) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8535)))) severity failure;
    assert RAM(8536) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8536)))) severity failure;
    assert RAM(8537) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8537)))) severity failure;
    assert RAM(8538) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8538)))) severity failure;
    assert RAM(8539) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8539)))) severity failure;
    assert RAM(8540) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8540)))) severity failure;
    assert RAM(8541) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8541)))) severity failure;
    assert RAM(8542) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8542)))) severity failure;
    assert RAM(8543) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8543)))) severity failure;
    assert RAM(8544) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8544)))) severity failure;
    assert RAM(8545) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8545)))) severity failure;
    assert RAM(8546) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8546)))) severity failure;
    assert RAM(8547) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8547)))) severity failure;
    assert RAM(8548) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8548)))) severity failure;
    assert RAM(8549) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8549)))) severity failure;
    assert RAM(8550) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8550)))) severity failure;
    assert RAM(8551) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8551)))) severity failure;
    assert RAM(8552) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8552)))) severity failure;
    assert RAM(8553) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8553)))) severity failure;
    assert RAM(8554) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8554)))) severity failure;
    assert RAM(8555) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8555)))) severity failure;
    assert RAM(8556) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8556)))) severity failure;
    assert RAM(8557) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8557)))) severity failure;
    assert RAM(8558) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8558)))) severity failure;
    assert RAM(8559) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8559)))) severity failure;
    assert RAM(8560) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8560)))) severity failure;
    assert RAM(8561) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8561)))) severity failure;
    assert RAM(8562) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8562)))) severity failure;
    assert RAM(8563) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8563)))) severity failure;
    assert RAM(8564) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8564)))) severity failure;
    assert RAM(8565) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8565)))) severity failure;
    assert RAM(8566) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8566)))) severity failure;
    assert RAM(8567) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8567)))) severity failure;
    assert RAM(8568) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8568)))) severity failure;
    assert RAM(8569) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8569)))) severity failure;
    assert RAM(8570) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8570)))) severity failure;
    assert RAM(8571) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8571)))) severity failure;
    assert RAM(8572) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8572)))) severity failure;
    assert RAM(8573) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8573)))) severity failure;
    assert RAM(8574) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8574)))) severity failure;
    assert RAM(8575) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8575)))) severity failure;
    assert RAM(8576) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8576)))) severity failure;
    assert RAM(8577) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8577)))) severity failure;
    assert RAM(8578) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8578)))) severity failure;
    assert RAM(8579) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8579)))) severity failure;
    assert RAM(8580) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8580)))) severity failure;
    assert RAM(8581) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8581)))) severity failure;
    assert RAM(8582) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8582)))) severity failure;
    assert RAM(8583) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8583)))) severity failure;
    assert RAM(8584) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8584)))) severity failure;
    assert RAM(8585) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8585)))) severity failure;
    assert RAM(8586) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8586)))) severity failure;
    assert RAM(8587) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8587)))) severity failure;
    assert RAM(8588) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8588)))) severity failure;
    assert RAM(8589) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8589)))) severity failure;
    assert RAM(8590) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8590)))) severity failure;
    assert RAM(8591) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8591)))) severity failure;
    assert RAM(8592) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8592)))) severity failure;
    assert RAM(8593) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8593)))) severity failure;
    assert RAM(8594) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8594)))) severity failure;
    assert RAM(8595) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8595)))) severity failure;
    assert RAM(8596) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8596)))) severity failure;
    assert RAM(8597) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8597)))) severity failure;
    assert RAM(8598) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8598)))) severity failure;
    assert RAM(8599) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8599)))) severity failure;
    assert RAM(8600) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8600)))) severity failure;
    assert RAM(8601) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8601)))) severity failure;
    assert RAM(8602) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8602)))) severity failure;
    assert RAM(8603) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8603)))) severity failure;
    assert RAM(8604) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8604)))) severity failure;
    assert RAM(8605) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8605)))) severity failure;
    assert RAM(8606) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8606)))) severity failure;
    assert RAM(8607) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8607)))) severity failure;
    assert RAM(8608) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8608)))) severity failure;
    assert RAM(8609) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8609)))) severity failure;
    assert RAM(8610) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8610)))) severity failure;
    assert RAM(8611) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8611)))) severity failure;
    assert RAM(8612) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8612)))) severity failure;
    assert RAM(8613) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8613)))) severity failure;
    assert RAM(8614) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8614)))) severity failure;
    assert RAM(8615) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8615)))) severity failure;
    assert RAM(8616) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8616)))) severity failure;
    assert RAM(8617) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8617)))) severity failure;
    assert RAM(8618) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8618)))) severity failure;
    assert RAM(8619) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8619)))) severity failure;
    assert RAM(8620) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8620)))) severity failure;
    assert RAM(8621) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8621)))) severity failure;
    assert RAM(8622) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8622)))) severity failure;
    assert RAM(8623) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8623)))) severity failure;
    assert RAM(8624) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8624)))) severity failure;
    assert RAM(8625) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8625)))) severity failure;
    assert RAM(8626) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8626)))) severity failure;
    assert RAM(8627) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8627)))) severity failure;
    assert RAM(8628) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8628)))) severity failure;
    assert RAM(8629) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8629)))) severity failure;
    assert RAM(8630) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8630)))) severity failure;
    assert RAM(8631) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8631)))) severity failure;
    assert RAM(8632) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8632)))) severity failure;
    assert RAM(8633) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8633)))) severity failure;
    assert RAM(8634) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8634)))) severity failure;
    assert RAM(8635) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8635)))) severity failure;
    assert RAM(8636) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8636)))) severity failure;
    assert RAM(8637) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8637)))) severity failure;
    assert RAM(8638) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8638)))) severity failure;
    assert RAM(8639) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8639)))) severity failure;
    assert RAM(8640) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8640)))) severity failure;
    assert RAM(8641) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8641)))) severity failure;
    assert RAM(8642) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8642)))) severity failure;
    assert RAM(8643) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8643)))) severity failure;
    assert RAM(8644) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8644)))) severity failure;
    assert RAM(8645) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8645)))) severity failure;
    assert RAM(8646) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8646)))) severity failure;
    assert RAM(8647) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8647)))) severity failure;
    assert RAM(8648) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8648)))) severity failure;
    assert RAM(8649) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8649)))) severity failure;
    assert RAM(8650) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8650)))) severity failure;
    assert RAM(8651) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8651)))) severity failure;
    assert RAM(8652) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8652)))) severity failure;
    assert RAM(8653) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8653)))) severity failure;
    assert RAM(8654) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8654)))) severity failure;
    assert RAM(8655) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8655)))) severity failure;
    assert RAM(8656) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8656)))) severity failure;
    assert RAM(8657) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8657)))) severity failure;
    assert RAM(8658) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8658)))) severity failure;
    assert RAM(8659) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8659)))) severity failure;
    assert RAM(8660) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8660)))) severity failure;
    assert RAM(8661) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8661)))) severity failure;
    assert RAM(8662) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8662)))) severity failure;
    assert RAM(8663) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8663)))) severity failure;
    assert RAM(8664) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8664)))) severity failure;
    assert RAM(8665) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8665)))) severity failure;
    assert RAM(8666) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8666)))) severity failure;
    assert RAM(8667) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8667)))) severity failure;
    assert RAM(8668) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8668)))) severity failure;
    assert RAM(8669) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8669)))) severity failure;
    assert RAM(8670) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8670)))) severity failure;
    assert RAM(8671) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8671)))) severity failure;
    assert RAM(8672) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8672)))) severity failure;
    assert RAM(8673) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8673)))) severity failure;
    assert RAM(8674) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8674)))) severity failure;
    assert RAM(8675) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8675)))) severity failure;
    assert RAM(8676) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8676)))) severity failure;
    assert RAM(8677) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8677)))) severity failure;
    assert RAM(8678) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8678)))) severity failure;
    assert RAM(8679) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8679)))) severity failure;
    assert RAM(8680) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8680)))) severity failure;
    assert RAM(8681) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8681)))) severity failure;
    assert RAM(8682) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8682)))) severity failure;
    assert RAM(8683) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8683)))) severity failure;
    assert RAM(8684) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8684)))) severity failure;
    assert RAM(8685) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8685)))) severity failure;
    assert RAM(8686) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8686)))) severity failure;
    assert RAM(8687) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8687)))) severity failure;
    assert RAM(8688) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8688)))) severity failure;
    assert RAM(8689) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8689)))) severity failure;
    assert RAM(8690) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8690)))) severity failure;
    assert RAM(8691) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8691)))) severity failure;
    assert RAM(8692) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8692)))) severity failure;
    assert RAM(8693) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8693)))) severity failure;
    assert RAM(8694) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8694)))) severity failure;
    assert RAM(8695) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8695)))) severity failure;
    assert RAM(8696) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8696)))) severity failure;
    assert RAM(8697) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8697)))) severity failure;
    assert RAM(8698) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8698)))) severity failure;
    assert RAM(8699) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8699)))) severity failure;
    assert RAM(8700) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8700)))) severity failure;
    assert RAM(8701) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8701)))) severity failure;
    assert RAM(8702) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8702)))) severity failure;
    assert RAM(8703) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8703)))) severity failure;
    assert RAM(8704) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8704)))) severity failure;
    assert RAM(8705) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8705)))) severity failure;
    assert RAM(8706) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8706)))) severity failure;
    assert RAM(8707) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8707)))) severity failure;
    assert RAM(8708) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8708)))) severity failure;
    assert RAM(8709) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8709)))) severity failure;
    assert RAM(8710) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8710)))) severity failure;
    assert RAM(8711) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8711)))) severity failure;
    assert RAM(8712) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8712)))) severity failure;
    assert RAM(8713) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8713)))) severity failure;
    assert RAM(8714) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8714)))) severity failure;
    assert RAM(8715) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8715)))) severity failure;
    assert RAM(8716) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8716)))) severity failure;
    assert RAM(8717) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8717)))) severity failure;
    assert RAM(8718) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8718)))) severity failure;
    assert RAM(8719) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8719)))) severity failure;
    assert RAM(8720) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8720)))) severity failure;
    assert RAM(8721) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8721)))) severity failure;
    assert RAM(8722) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8722)))) severity failure;
    assert RAM(8723) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8723)))) severity failure;
    assert RAM(8724) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8724)))) severity failure;
    assert RAM(8725) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8725)))) severity failure;
    assert RAM(8726) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8726)))) severity failure;
    assert RAM(8727) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8727)))) severity failure;
    assert RAM(8728) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8728)))) severity failure;
    assert RAM(8729) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8729)))) severity failure;
    assert RAM(8730) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8730)))) severity failure;
    assert RAM(8731) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8731)))) severity failure;
    assert RAM(8732) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8732)))) severity failure;
    assert RAM(8733) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8733)))) severity failure;
    assert RAM(8734) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8734)))) severity failure;
    assert RAM(8735) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8735)))) severity failure;
    assert RAM(8736) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8736)))) severity failure;
    assert RAM(8737) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8737)))) severity failure;
    assert RAM(8738) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8738)))) severity failure;
    assert RAM(8739) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8739)))) severity failure;
    assert RAM(8740) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8740)))) severity failure;
    assert RAM(8741) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8741)))) severity failure;
    assert RAM(8742) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8742)))) severity failure;
    assert RAM(8743) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8743)))) severity failure;
    assert RAM(8744) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8744)))) severity failure;
    assert RAM(8745) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8745)))) severity failure;
    assert RAM(8746) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8746)))) severity failure;
    assert RAM(8747) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8747)))) severity failure;
    assert RAM(8748) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8748)))) severity failure;
    assert RAM(8749) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8749)))) severity failure;
    assert RAM(8750) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8750)))) severity failure;
    assert RAM(8751) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8751)))) severity failure;
    assert RAM(8752) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8752)))) severity failure;
    assert RAM(8753) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8753)))) severity failure;
    assert RAM(8754) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8754)))) severity failure;
    assert RAM(8755) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8755)))) severity failure;
    assert RAM(8756) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8756)))) severity failure;
    assert RAM(8757) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8757)))) severity failure;
    assert RAM(8758) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8758)))) severity failure;
    assert RAM(8759) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8759)))) severity failure;
    assert RAM(8760) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8760)))) severity failure;
    assert RAM(8761) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8761)))) severity failure;
    assert RAM(8762) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8762)))) severity failure;
    assert RAM(8763) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8763)))) severity failure;
    assert RAM(8764) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8764)))) severity failure;
    assert RAM(8765) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8765)))) severity failure;
    assert RAM(8766) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8766)))) severity failure;
    assert RAM(8767) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8767)))) severity failure;
    assert RAM(8768) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8768)))) severity failure;
    assert RAM(8769) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8769)))) severity failure;
    assert RAM(8770) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8770)))) severity failure;
    assert RAM(8771) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8771)))) severity failure;
    assert RAM(8772) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8772)))) severity failure;
    assert RAM(8773) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8773)))) severity failure;
    assert RAM(8774) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8774)))) severity failure;
    assert RAM(8775) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8775)))) severity failure;
    assert RAM(8776) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8776)))) severity failure;
    assert RAM(8777) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8777)))) severity failure;
    assert RAM(8778) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8778)))) severity failure;
    assert RAM(8779) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8779)))) severity failure;
    assert RAM(8780) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8780)))) severity failure;
    assert RAM(8781) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8781)))) severity failure;
    assert RAM(8782) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8782)))) severity failure;
    assert RAM(8783) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8783)))) severity failure;
    assert RAM(8784) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8784)))) severity failure;
    assert RAM(8785) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8785)))) severity failure;
    assert RAM(8786) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8786)))) severity failure;
    assert RAM(8787) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8787)))) severity failure;
    assert RAM(8788) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8788)))) severity failure;
    assert RAM(8789) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8789)))) severity failure;
    assert RAM(8790) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8790)))) severity failure;
    assert RAM(8791) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8791)))) severity failure;
    assert RAM(8792) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8792)))) severity failure;
    assert RAM(8793) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8793)))) severity failure;
    assert RAM(8794) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8794)))) severity failure;
    assert RAM(8795) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8795)))) severity failure;
    assert RAM(8796) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8796)))) severity failure;
    assert RAM(8797) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8797)))) severity failure;
    assert RAM(8798) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8798)))) severity failure;
    assert RAM(8799) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8799)))) severity failure;
    assert RAM(8800) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8800)))) severity failure;
    assert RAM(8801) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8801)))) severity failure;
    assert RAM(8802) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8802)))) severity failure;
    assert RAM(8803) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8803)))) severity failure;
    assert RAM(8804) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8804)))) severity failure;
    assert RAM(8805) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8805)))) severity failure;
    assert RAM(8806) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8806)))) severity failure;
    assert RAM(8807) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8807)))) severity failure;
    assert RAM(8808) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8808)))) severity failure;
    assert RAM(8809) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8809)))) severity failure;
    assert RAM(8810) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8810)))) severity failure;
    assert RAM(8811) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8811)))) severity failure;
    assert RAM(8812) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8812)))) severity failure;
    assert RAM(8813) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8813)))) severity failure;
    assert RAM(8814) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8814)))) severity failure;
    assert RAM(8815) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8815)))) severity failure;
    assert RAM(8816) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8816)))) severity failure;
    assert RAM(8817) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8817)))) severity failure;
    assert RAM(8818) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8818)))) severity failure;
    assert RAM(8819) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8819)))) severity failure;
    assert RAM(8820) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8820)))) severity failure;
    assert RAM(8821) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8821)))) severity failure;
    assert RAM(8822) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8822)))) severity failure;
    assert RAM(8823) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8823)))) severity failure;
    assert RAM(8824) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8824)))) severity failure;
    assert RAM(8825) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8825)))) severity failure;
    assert RAM(8826) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8826)))) severity failure;
    assert RAM(8827) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8827)))) severity failure;
    assert RAM(8828) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8828)))) severity failure;
    assert RAM(8829) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8829)))) severity failure;
    assert RAM(8830) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8830)))) severity failure;
    assert RAM(8831) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8831)))) severity failure;
    assert RAM(8832) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8832)))) severity failure;
    assert RAM(8833) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8833)))) severity failure;
    assert RAM(8834) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8834)))) severity failure;
    assert RAM(8835) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8835)))) severity failure;
    assert RAM(8836) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8836)))) severity failure;
    assert RAM(8837) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8837)))) severity failure;
    assert RAM(8838) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8838)))) severity failure;
    assert RAM(8839) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8839)))) severity failure;
    assert RAM(8840) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8840)))) severity failure;
    assert RAM(8841) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8841)))) severity failure;
    assert RAM(8842) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8842)))) severity failure;
    assert RAM(8843) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8843)))) severity failure;
    assert RAM(8844) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8844)))) severity failure;
    assert RAM(8845) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8845)))) severity failure;
    assert RAM(8846) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8846)))) severity failure;
    assert RAM(8847) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8847)))) severity failure;
    assert RAM(8848) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8848)))) severity failure;
    assert RAM(8849) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8849)))) severity failure;
    assert RAM(8850) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8850)))) severity failure;
    assert RAM(8851) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8851)))) severity failure;
    assert RAM(8852) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8852)))) severity failure;
    assert RAM(8853) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8853)))) severity failure;
    assert RAM(8854) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8854)))) severity failure;
    assert RAM(8855) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8855)))) severity failure;
    assert RAM(8856) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8856)))) severity failure;
    assert RAM(8857) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8857)))) severity failure;
    assert RAM(8858) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8858)))) severity failure;
    assert RAM(8859) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8859)))) severity failure;
    assert RAM(8860) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8860)))) severity failure;
    assert RAM(8861) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8861)))) severity failure;
    assert RAM(8862) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8862)))) severity failure;
    assert RAM(8863) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8863)))) severity failure;
    assert RAM(8864) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8864)))) severity failure;
    assert RAM(8865) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8865)))) severity failure;
    assert RAM(8866) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8866)))) severity failure;
    assert RAM(8867) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8867)))) severity failure;
    assert RAM(8868) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8868)))) severity failure;
    assert RAM(8869) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8869)))) severity failure;
    assert RAM(8870) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8870)))) severity failure;
    assert RAM(8871) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8871)))) severity failure;
    assert RAM(8872) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8872)))) severity failure;
    assert RAM(8873) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8873)))) severity failure;
    assert RAM(8874) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8874)))) severity failure;
    assert RAM(8875) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8875)))) severity failure;
    assert RAM(8876) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8876)))) severity failure;
    assert RAM(8877) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8877)))) severity failure;
    assert RAM(8878) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8878)))) severity failure;
    assert RAM(8879) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8879)))) severity failure;
    assert RAM(8880) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8880)))) severity failure;
    assert RAM(8881) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8881)))) severity failure;
    assert RAM(8882) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8882)))) severity failure;
    assert RAM(8883) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8883)))) severity failure;
    assert RAM(8884) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8884)))) severity failure;
    assert RAM(8885) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8885)))) severity failure;
    assert RAM(8886) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8886)))) severity failure;
    assert RAM(8887) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8887)))) severity failure;
    assert RAM(8888) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8888)))) severity failure;
    assert RAM(8889) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8889)))) severity failure;
    assert RAM(8890) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8890)))) severity failure;
    assert RAM(8891) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8891)))) severity failure;
    assert RAM(8892) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8892)))) severity failure;
    assert RAM(8893) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8893)))) severity failure;
    assert RAM(8894) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8894)))) severity failure;
    assert RAM(8895) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8895)))) severity failure;
    assert RAM(8896) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8896)))) severity failure;
    assert RAM(8897) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8897)))) severity failure;
    assert RAM(8898) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8898)))) severity failure;
    assert RAM(8899) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8899)))) severity failure;
    assert RAM(8900) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8900)))) severity failure;
    assert RAM(8901) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8901)))) severity failure;
    assert RAM(8902) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8902)))) severity failure;
    assert RAM(8903) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8903)))) severity failure;
    assert RAM(8904) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8904)))) severity failure;
    assert RAM(8905) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8905)))) severity failure;
    assert RAM(8906) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8906)))) severity failure;
    assert RAM(8907) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8907)))) severity failure;
    assert RAM(8908) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8908)))) severity failure;
    assert RAM(8909) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8909)))) severity failure;
    assert RAM(8910) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8910)))) severity failure;
    assert RAM(8911) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8911)))) severity failure;
    assert RAM(8912) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8912)))) severity failure;
    assert RAM(8913) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8913)))) severity failure;
    assert RAM(8914) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8914)))) severity failure;
    assert RAM(8915) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8915)))) severity failure;
    assert RAM(8916) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8916)))) severity failure;
    assert RAM(8917) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8917)))) severity failure;
    assert RAM(8918) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8918)))) severity failure;
    assert RAM(8919) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8919)))) severity failure;
    assert RAM(8920) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8920)))) severity failure;
    assert RAM(8921) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8921)))) severity failure;
    assert RAM(8922) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8922)))) severity failure;
    assert RAM(8923) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8923)))) severity failure;
    assert RAM(8924) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8924)))) severity failure;
    assert RAM(8925) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8925)))) severity failure;
    assert RAM(8926) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8926)))) severity failure;
    assert RAM(8927) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8927)))) severity failure;
    assert RAM(8928) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8928)))) severity failure;
    assert RAM(8929) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8929)))) severity failure;
    assert RAM(8930) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8930)))) severity failure;
    assert RAM(8931) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8931)))) severity failure;
    assert RAM(8932) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8932)))) severity failure;
    assert RAM(8933) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8933)))) severity failure;
    assert RAM(8934) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8934)))) severity failure;
    assert RAM(8935) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8935)))) severity failure;
    assert RAM(8936) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8936)))) severity failure;
    assert RAM(8937) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8937)))) severity failure;
    assert RAM(8938) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8938)))) severity failure;
    assert RAM(8939) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8939)))) severity failure;
    assert RAM(8940) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8940)))) severity failure;
    assert RAM(8941) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8941)))) severity failure;
    assert RAM(8942) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8942)))) severity failure;
    assert RAM(8943) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8943)))) severity failure;
    assert RAM(8944) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8944)))) severity failure;
    assert RAM(8945) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8945)))) severity failure;
    assert RAM(8946) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8946)))) severity failure;
    assert RAM(8947) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8947)))) severity failure;
    assert RAM(8948) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8948)))) severity failure;
    assert RAM(8949) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8949)))) severity failure;
    assert RAM(8950) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8950)))) severity failure;
    assert RAM(8951) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8951)))) severity failure;
    assert RAM(8952) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8952)))) severity failure;
    assert RAM(8953) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8953)))) severity failure;
    assert RAM(8954) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8954)))) severity failure;
    assert RAM(8955) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8955)))) severity failure;
    assert RAM(8956) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8956)))) severity failure;
    assert RAM(8957) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8957)))) severity failure;
    assert RAM(8958) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8958)))) severity failure;
    assert RAM(8959) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8959)))) severity failure;
    assert RAM(8960) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8960)))) severity failure;
    assert RAM(8961) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8961)))) severity failure;
    assert RAM(8962) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8962)))) severity failure;
    assert RAM(8963) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8963)))) severity failure;
    assert RAM(8964) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8964)))) severity failure;
    assert RAM(8965) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8965)))) severity failure;
    assert RAM(8966) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8966)))) severity failure;
    assert RAM(8967) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8967)))) severity failure;
    assert RAM(8968) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8968)))) severity failure;
    assert RAM(8969) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8969)))) severity failure;
    assert RAM(8970) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8970)))) severity failure;
    assert RAM(8971) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8971)))) severity failure;
    assert RAM(8972) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8972)))) severity failure;
    assert RAM(8973) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8973)))) severity failure;
    assert RAM(8974) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8974)))) severity failure;
    assert RAM(8975) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8975)))) severity failure;
    assert RAM(8976) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8976)))) severity failure;
    assert RAM(8977) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8977)))) severity failure;
    assert RAM(8978) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8978)))) severity failure;
    assert RAM(8979) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8979)))) severity failure;
    assert RAM(8980) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8980)))) severity failure;
    assert RAM(8981) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8981)))) severity failure;
    assert RAM(8982) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8982)))) severity failure;
    assert RAM(8983) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8983)))) severity failure;
    assert RAM(8984) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8984)))) severity failure;
    assert RAM(8985) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8985)))) severity failure;
    assert RAM(8986) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8986)))) severity failure;
    assert RAM(8987) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8987)))) severity failure;
    assert RAM(8988) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8988)))) severity failure;
    assert RAM(8989) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8989)))) severity failure;
    assert RAM(8990) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8990)))) severity failure;
    assert RAM(8991) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8991)))) severity failure;
    assert RAM(8992) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8992)))) severity failure;
    assert RAM(8993) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8993)))) severity failure;
    assert RAM(8994) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8994)))) severity failure;
    assert RAM(8995) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8995)))) severity failure;
    assert RAM(8996) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8996)))) severity failure;
    assert RAM(8997) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8997)))) severity failure;
    assert RAM(8998) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(8998)))) severity failure;
    assert RAM(8999) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(8999)))) severity failure;
    assert RAM(9000) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9000)))) severity failure;
    assert RAM(9001) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9001)))) severity failure;
    assert RAM(9002) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9002)))) severity failure;
    assert RAM(9003) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9003)))) severity failure;
    assert RAM(9004) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9004)))) severity failure;
    assert RAM(9005) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9005)))) severity failure;
    assert RAM(9006) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9006)))) severity failure;
    assert RAM(9007) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9007)))) severity failure;
    assert RAM(9008) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9008)))) severity failure;
    assert RAM(9009) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9009)))) severity failure;
    assert RAM(9010) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9010)))) severity failure;
    assert RAM(9011) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9011)))) severity failure;
    assert RAM(9012) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9012)))) severity failure;
    assert RAM(9013) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9013)))) severity failure;
    assert RAM(9014) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9014)))) severity failure;
    assert RAM(9015) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9015)))) severity failure;
    assert RAM(9016) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9016)))) severity failure;
    assert RAM(9017) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9017)))) severity failure;
    assert RAM(9018) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9018)))) severity failure;
    assert RAM(9019) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9019)))) severity failure;
    assert RAM(9020) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9020)))) severity failure;
    assert RAM(9021) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9021)))) severity failure;
    assert RAM(9022) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9022)))) severity failure;
    assert RAM(9023) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9023)))) severity failure;
    assert RAM(9024) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9024)))) severity failure;
    assert RAM(9025) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9025)))) severity failure;
    assert RAM(9026) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9026)))) severity failure;
    assert RAM(9027) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9027)))) severity failure;
    assert RAM(9028) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9028)))) severity failure;
    assert RAM(9029) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9029)))) severity failure;
    assert RAM(9030) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9030)))) severity failure;
    assert RAM(9031) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9031)))) severity failure;
    assert RAM(9032) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9032)))) severity failure;
    assert RAM(9033) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9033)))) severity failure;
    assert RAM(9034) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9034)))) severity failure;
    assert RAM(9035) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9035)))) severity failure;
    assert RAM(9036) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9036)))) severity failure;
    assert RAM(9037) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9037)))) severity failure;
    assert RAM(9038) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9038)))) severity failure;
    assert RAM(9039) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9039)))) severity failure;
    assert RAM(9040) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9040)))) severity failure;
    assert RAM(9041) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9041)))) severity failure;
    assert RAM(9042) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9042)))) severity failure;
    assert RAM(9043) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9043)))) severity failure;
    assert RAM(9044) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9044)))) severity failure;
    assert RAM(9045) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9045)))) severity failure;
    assert RAM(9046) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9046)))) severity failure;
    assert RAM(9047) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9047)))) severity failure;
    assert RAM(9048) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9048)))) severity failure;
    assert RAM(9049) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9049)))) severity failure;
    assert RAM(9050) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9050)))) severity failure;
    assert RAM(9051) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9051)))) severity failure;
    assert RAM(9052) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9052)))) severity failure;
    assert RAM(9053) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9053)))) severity failure;
    assert RAM(9054) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9054)))) severity failure;
    assert RAM(9055) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9055)))) severity failure;
    assert RAM(9056) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9056)))) severity failure;
    assert RAM(9057) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9057)))) severity failure;
    assert RAM(9058) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9058)))) severity failure;
    assert RAM(9059) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9059)))) severity failure;
    assert RAM(9060) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9060)))) severity failure;
    assert RAM(9061) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9061)))) severity failure;
    assert RAM(9062) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9062)))) severity failure;
    assert RAM(9063) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9063)))) severity failure;
    assert RAM(9064) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9064)))) severity failure;
    assert RAM(9065) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9065)))) severity failure;
    assert RAM(9066) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9066)))) severity failure;
    assert RAM(9067) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9067)))) severity failure;
    assert RAM(9068) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9068)))) severity failure;
    assert RAM(9069) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9069)))) severity failure;
    assert RAM(9070) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9070)))) severity failure;
    assert RAM(9071) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9071)))) severity failure;
    assert RAM(9072) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9072)))) severity failure;
    assert RAM(9073) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9073)))) severity failure;
    assert RAM(9074) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9074)))) severity failure;
    assert RAM(9075) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9075)))) severity failure;
    assert RAM(9076) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9076)))) severity failure;
    assert RAM(9077) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9077)))) severity failure;
    assert RAM(9078) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9078)))) severity failure;
    assert RAM(9079) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9079)))) severity failure;
    assert RAM(9080) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9080)))) severity failure;
    assert RAM(9081) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9081)))) severity failure;
    assert RAM(9082) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9082)))) severity failure;
    assert RAM(9083) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9083)))) severity failure;
    assert RAM(9084) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9084)))) severity failure;
    assert RAM(9085) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9085)))) severity failure;
    assert RAM(9086) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9086)))) severity failure;
    assert RAM(9087) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9087)))) severity failure;
    assert RAM(9088) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9088)))) severity failure;
    assert RAM(9089) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9089)))) severity failure;
    assert RAM(9090) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9090)))) severity failure;
    assert RAM(9091) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9091)))) severity failure;
    assert RAM(9092) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9092)))) severity failure;
    assert RAM(9093) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9093)))) severity failure;
    assert RAM(9094) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9094)))) severity failure;
    assert RAM(9095) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9095)))) severity failure;
    assert RAM(9096) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9096)))) severity failure;
    assert RAM(9097) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9097)))) severity failure;
    assert RAM(9098) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9098)))) severity failure;
    assert RAM(9099) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9099)))) severity failure;
    assert RAM(9100) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9100)))) severity failure;
    assert RAM(9101) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9101)))) severity failure;
    assert RAM(9102) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9102)))) severity failure;
    assert RAM(9103) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9103)))) severity failure;
    assert RAM(9104) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9104)))) severity failure;
    assert RAM(9105) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9105)))) severity failure;
    assert RAM(9106) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9106)))) severity failure;
    assert RAM(9107) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9107)))) severity failure;
    assert RAM(9108) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9108)))) severity failure;
    assert RAM(9109) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9109)))) severity failure;
    assert RAM(9110) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9110)))) severity failure;
    assert RAM(9111) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9111)))) severity failure;
    assert RAM(9112) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9112)))) severity failure;
    assert RAM(9113) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9113)))) severity failure;
    assert RAM(9114) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9114)))) severity failure;
    assert RAM(9115) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9115)))) severity failure;
    assert RAM(9116) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9116)))) severity failure;
    assert RAM(9117) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9117)))) severity failure;
    assert RAM(9118) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9118)))) severity failure;
    assert RAM(9119) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9119)))) severity failure;
    assert RAM(9120) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9120)))) severity failure;
    assert RAM(9121) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9121)))) severity failure;
    assert RAM(9122) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9122)))) severity failure;
    assert RAM(9123) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9123)))) severity failure;
    assert RAM(9124) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9124)))) severity failure;
    assert RAM(9125) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9125)))) severity failure;
    assert RAM(9126) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9126)))) severity failure;
    assert RAM(9127) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9127)))) severity failure;
    assert RAM(9128) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9128)))) severity failure;
    assert RAM(9129) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9129)))) severity failure;
    assert RAM(9130) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9130)))) severity failure;
    assert RAM(9131) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9131)))) severity failure;
    assert RAM(9132) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9132)))) severity failure;
    assert RAM(9133) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9133)))) severity failure;
    assert RAM(9134) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9134)))) severity failure;
    assert RAM(9135) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9135)))) severity failure;
    assert RAM(9136) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9136)))) severity failure;
    assert RAM(9137) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9137)))) severity failure;
    assert RAM(9138) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9138)))) severity failure;
    assert RAM(9139) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9139)))) severity failure;
    assert RAM(9140) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9140)))) severity failure;
    assert RAM(9141) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9141)))) severity failure;
    assert RAM(9142) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9142)))) severity failure;
    assert RAM(9143) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9143)))) severity failure;
    assert RAM(9144) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9144)))) severity failure;
    assert RAM(9145) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9145)))) severity failure;
    assert RAM(9146) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9146)))) severity failure;
    assert RAM(9147) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9147)))) severity failure;
    assert RAM(9148) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9148)))) severity failure;
    assert RAM(9149) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9149)))) severity failure;
    assert RAM(9150) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9150)))) severity failure;
    assert RAM(9151) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9151)))) severity failure;
    assert RAM(9152) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9152)))) severity failure;
    assert RAM(9153) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9153)))) severity failure;
    assert RAM(9154) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9154)))) severity failure;
    assert RAM(9155) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9155)))) severity failure;
    assert RAM(9156) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9156)))) severity failure;
    assert RAM(9157) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9157)))) severity failure;
    assert RAM(9158) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9158)))) severity failure;
    assert RAM(9159) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9159)))) severity failure;
    assert RAM(9160) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9160)))) severity failure;
    assert RAM(9161) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9161)))) severity failure;
    assert RAM(9162) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9162)))) severity failure;
    assert RAM(9163) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9163)))) severity failure;
    assert RAM(9164) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9164)))) severity failure;
    assert RAM(9165) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9165)))) severity failure;
    assert RAM(9166) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9166)))) severity failure;
    assert RAM(9167) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9167)))) severity failure;
    assert RAM(9168) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9168)))) severity failure;
    assert RAM(9169) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9169)))) severity failure;
    assert RAM(9170) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9170)))) severity failure;
    assert RAM(9171) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9171)))) severity failure;
    assert RAM(9172) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9172)))) severity failure;
    assert RAM(9173) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9173)))) severity failure;
    assert RAM(9174) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9174)))) severity failure;
    assert RAM(9175) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9175)))) severity failure;
    assert RAM(9176) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9176)))) severity failure;
    assert RAM(9177) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9177)))) severity failure;
    assert RAM(9178) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9178)))) severity failure;
    assert RAM(9179) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9179)))) severity failure;
    assert RAM(9180) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9180)))) severity failure;
    assert RAM(9181) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9181)))) severity failure;
    assert RAM(9182) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9182)))) severity failure;
    assert RAM(9183) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9183)))) severity failure;
    assert RAM(9184) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9184)))) severity failure;
    assert RAM(9185) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9185)))) severity failure;
    assert RAM(9186) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9186)))) severity failure;
    assert RAM(9187) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9187)))) severity failure;
    assert RAM(9188) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9188)))) severity failure;
    assert RAM(9189) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9189)))) severity failure;
    assert RAM(9190) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9190)))) severity failure;
    assert RAM(9191) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9191)))) severity failure;
    assert RAM(9192) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9192)))) severity failure;
    assert RAM(9193) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9193)))) severity failure;
    assert RAM(9194) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9194)))) severity failure;
    assert RAM(9195) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9195)))) severity failure;
    assert RAM(9196) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9196)))) severity failure;
    assert RAM(9197) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9197)))) severity failure;
    assert RAM(9198) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9198)))) severity failure;
    assert RAM(9199) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9199)))) severity failure;
    assert RAM(9200) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9200)))) severity failure;
    assert RAM(9201) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9201)))) severity failure;
    assert RAM(9202) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9202)))) severity failure;
    assert RAM(9203) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9203)))) severity failure;
    assert RAM(9204) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9204)))) severity failure;
    assert RAM(9205) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9205)))) severity failure;
    assert RAM(9206) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9206)))) severity failure;
    assert RAM(9207) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9207)))) severity failure;
    assert RAM(9208) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9208)))) severity failure;
    assert RAM(9209) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9209)))) severity failure;
    assert RAM(9210) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9210)))) severity failure;
    assert RAM(9211) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9211)))) severity failure;
    assert RAM(9212) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9212)))) severity failure;
    assert RAM(9213) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9213)))) severity failure;
    assert RAM(9214) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9214)))) severity failure;
    assert RAM(9215) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9215)))) severity failure;
    assert RAM(9216) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9216)))) severity failure;
    assert RAM(9217) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9217)))) severity failure;
    assert RAM(9218) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9218)))) severity failure;
    assert RAM(9219) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9219)))) severity failure;
    assert RAM(9220) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9220)))) severity failure;
    assert RAM(9221) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9221)))) severity failure;
    assert RAM(9222) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9222)))) severity failure;
    assert RAM(9223) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9223)))) severity failure;
    assert RAM(9224) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9224)))) severity failure;
    assert RAM(9225) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9225)))) severity failure;
    assert RAM(9226) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9226)))) severity failure;
    assert RAM(9227) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9227)))) severity failure;
    assert RAM(9228) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9228)))) severity failure;
    assert RAM(9229) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9229)))) severity failure;
    assert RAM(9230) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9230)))) severity failure;
    assert RAM(9231) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9231)))) severity failure;
    assert RAM(9232) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9232)))) severity failure;
    assert RAM(9233) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9233)))) severity failure;
    assert RAM(9234) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9234)))) severity failure;
    assert RAM(9235) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9235)))) severity failure;
    assert RAM(9236) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9236)))) severity failure;
    assert RAM(9237) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9237)))) severity failure;
    assert RAM(9238) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9238)))) severity failure;
    assert RAM(9239) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9239)))) severity failure;
    assert RAM(9240) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9240)))) severity failure;
    assert RAM(9241) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9241)))) severity failure;
    assert RAM(9242) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9242)))) severity failure;
    assert RAM(9243) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9243)))) severity failure;
    assert RAM(9244) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9244)))) severity failure;
    assert RAM(9245) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9245)))) severity failure;
    assert RAM(9246) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9246)))) severity failure;
    assert RAM(9247) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9247)))) severity failure;
    assert RAM(9248) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9248)))) severity failure;
    assert RAM(9249) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9249)))) severity failure;
    assert RAM(9250) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9250)))) severity failure;
    assert RAM(9251) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9251)))) severity failure;
    assert RAM(9252) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9252)))) severity failure;
    assert RAM(9253) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9253)))) severity failure;
    assert RAM(9254) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9254)))) severity failure;
    assert RAM(9255) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9255)))) severity failure;
    assert RAM(9256) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9256)))) severity failure;
    assert RAM(9257) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9257)))) severity failure;
    assert RAM(9258) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9258)))) severity failure;
    assert RAM(9259) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9259)))) severity failure;
    assert RAM(9260) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9260)))) severity failure;
    assert RAM(9261) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9261)))) severity failure;
    assert RAM(9262) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9262)))) severity failure;
    assert RAM(9263) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9263)))) severity failure;
    assert RAM(9264) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9264)))) severity failure;
    assert RAM(9265) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9265)))) severity failure;
    assert RAM(9266) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9266)))) severity failure;
    assert RAM(9267) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9267)))) severity failure;
    assert RAM(9268) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9268)))) severity failure;
    assert RAM(9269) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9269)))) severity failure;
    assert RAM(9270) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9270)))) severity failure;
    assert RAM(9271) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9271)))) severity failure;
    assert RAM(9272) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9272)))) severity failure;
    assert RAM(9273) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9273)))) severity failure;
    assert RAM(9274) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9274)))) severity failure;
    assert RAM(9275) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9275)))) severity failure;
    assert RAM(9276) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9276)))) severity failure;
    assert RAM(9277) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9277)))) severity failure;
    assert RAM(9278) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9278)))) severity failure;
    assert RAM(9279) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9279)))) severity failure;
    assert RAM(9280) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9280)))) severity failure;
    assert RAM(9281) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9281)))) severity failure;
    assert RAM(9282) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9282)))) severity failure;
    assert RAM(9283) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9283)))) severity failure;
    assert RAM(9284) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9284)))) severity failure;
    assert RAM(9285) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9285)))) severity failure;
    assert RAM(9286) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9286)))) severity failure;
    assert RAM(9287) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9287)))) severity failure;
    assert RAM(9288) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9288)))) severity failure;
    assert RAM(9289) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9289)))) severity failure;
    assert RAM(9290) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9290)))) severity failure;
    assert RAM(9291) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9291)))) severity failure;
    assert RAM(9292) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9292)))) severity failure;
    assert RAM(9293) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9293)))) severity failure;
    assert RAM(9294) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9294)))) severity failure;
    assert RAM(9295) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9295)))) severity failure;
    assert RAM(9296) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9296)))) severity failure;
    assert RAM(9297) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9297)))) severity failure;
    assert RAM(9298) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9298)))) severity failure;
    assert RAM(9299) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9299)))) severity failure;
    assert RAM(9300) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9300)))) severity failure;
    assert RAM(9301) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9301)))) severity failure;
    assert RAM(9302) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9302)))) severity failure;
    assert RAM(9303) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9303)))) severity failure;
    assert RAM(9304) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9304)))) severity failure;
    assert RAM(9305) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9305)))) severity failure;
    assert RAM(9306) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9306)))) severity failure;
    assert RAM(9307) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9307)))) severity failure;
    assert RAM(9308) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9308)))) severity failure;
    assert RAM(9309) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9309)))) severity failure;
    assert RAM(9310) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9310)))) severity failure;
    assert RAM(9311) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9311)))) severity failure;
    assert RAM(9312) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9312)))) severity failure;
    assert RAM(9313) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9313)))) severity failure;
    assert RAM(9314) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9314)))) severity failure;
    assert RAM(9315) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9315)))) severity failure;
    assert RAM(9316) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9316)))) severity failure;
    assert RAM(9317) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9317)))) severity failure;
    assert RAM(9318) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9318)))) severity failure;
    assert RAM(9319) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9319)))) severity failure;
    assert RAM(9320) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9320)))) severity failure;
    assert RAM(9321) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9321)))) severity failure;
    assert RAM(9322) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9322)))) severity failure;
    assert RAM(9323) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9323)))) severity failure;
    assert RAM(9324) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9324)))) severity failure;
    assert RAM(9325) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9325)))) severity failure;
    assert RAM(9326) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9326)))) severity failure;
    assert RAM(9327) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9327)))) severity failure;
    assert RAM(9328) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9328)))) severity failure;
    assert RAM(9329) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9329)))) severity failure;
    assert RAM(9330) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9330)))) severity failure;
    assert RAM(9331) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9331)))) severity failure;
    assert RAM(9332) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9332)))) severity failure;
    assert RAM(9333) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9333)))) severity failure;
    assert RAM(9334) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9334)))) severity failure;
    assert RAM(9335) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9335)))) severity failure;
    assert RAM(9336) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9336)))) severity failure;
    assert RAM(9337) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9337)))) severity failure;
    assert RAM(9338) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9338)))) severity failure;
    assert RAM(9339) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9339)))) severity failure;
    assert RAM(9340) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9340)))) severity failure;
    assert RAM(9341) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9341)))) severity failure;
    assert RAM(9342) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9342)))) severity failure;
    assert RAM(9343) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9343)))) severity failure;
    assert RAM(9344) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9344)))) severity failure;
    assert RAM(9345) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9345)))) severity failure;
    assert RAM(9346) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9346)))) severity failure;
    assert RAM(9347) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9347)))) severity failure;
    assert RAM(9348) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9348)))) severity failure;
    assert RAM(9349) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9349)))) severity failure;
    assert RAM(9350) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9350)))) severity failure;
    assert RAM(9351) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9351)))) severity failure;
    assert RAM(9352) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9352)))) severity failure;
    assert RAM(9353) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9353)))) severity failure;
    assert RAM(9354) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9354)))) severity failure;
    assert RAM(9355) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9355)))) severity failure;
    assert RAM(9356) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9356)))) severity failure;
    assert RAM(9357) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9357)))) severity failure;
    assert RAM(9358) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9358)))) severity failure;
    assert RAM(9359) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9359)))) severity failure;
    assert RAM(9360) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9360)))) severity failure;
    assert RAM(9361) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9361)))) severity failure;
    assert RAM(9362) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9362)))) severity failure;
    assert RAM(9363) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9363)))) severity failure;
    assert RAM(9364) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9364)))) severity failure;
    assert RAM(9365) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9365)))) severity failure;
    assert RAM(9366) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9366)))) severity failure;
    assert RAM(9367) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9367)))) severity failure;
    assert RAM(9368) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9368)))) severity failure;
    assert RAM(9369) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9369)))) severity failure;
    assert RAM(9370) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9370)))) severity failure;
    assert RAM(9371) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9371)))) severity failure;
    assert RAM(9372) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9372)))) severity failure;
    assert RAM(9373) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9373)))) severity failure;
    assert RAM(9374) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9374)))) severity failure;
    assert RAM(9375) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9375)))) severity failure;
    assert RAM(9376) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9376)))) severity failure;
    assert RAM(9377) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9377)))) severity failure;
    assert RAM(9378) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9378)))) severity failure;
    assert RAM(9379) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9379)))) severity failure;
    assert RAM(9380) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9380)))) severity failure;
    assert RAM(9381) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9381)))) severity failure;
    assert RAM(9382) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9382)))) severity failure;
    assert RAM(9383) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9383)))) severity failure;
    assert RAM(9384) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9384)))) severity failure;
    assert RAM(9385) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9385)))) severity failure;
    assert RAM(9386) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9386)))) severity failure;
    assert RAM(9387) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9387)))) severity failure;
    assert RAM(9388) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9388)))) severity failure;
    assert RAM(9389) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9389)))) severity failure;
    assert RAM(9390) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9390)))) severity failure;
    assert RAM(9391) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9391)))) severity failure;
    assert RAM(9392) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9392)))) severity failure;
    assert RAM(9393) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9393)))) severity failure;
    assert RAM(9394) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9394)))) severity failure;
    assert RAM(9395) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9395)))) severity failure;
    assert RAM(9396) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9396)))) severity failure;
    assert RAM(9397) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9397)))) severity failure;
    assert RAM(9398) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9398)))) severity failure;
    assert RAM(9399) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9399)))) severity failure;
    assert RAM(9400) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9400)))) severity failure;
    assert RAM(9401) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9401)))) severity failure;
    assert RAM(9402) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9402)))) severity failure;
    assert RAM(9403) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9403)))) severity failure;
    assert RAM(9404) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9404)))) severity failure;
    assert RAM(9405) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9405)))) severity failure;
    assert RAM(9406) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9406)))) severity failure;
    assert RAM(9407) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9407)))) severity failure;
    assert RAM(9408) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9408)))) severity failure;
    assert RAM(9409) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9409)))) severity failure;
    assert RAM(9410) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9410)))) severity failure;
    assert RAM(9411) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9411)))) severity failure;
    assert RAM(9412) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9412)))) severity failure;
    assert RAM(9413) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9413)))) severity failure;
    assert RAM(9414) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9414)))) severity failure;
    assert RAM(9415) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9415)))) severity failure;
    assert RAM(9416) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9416)))) severity failure;
    assert RAM(9417) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9417)))) severity failure;
    assert RAM(9418) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9418)))) severity failure;
    assert RAM(9419) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9419)))) severity failure;
    assert RAM(9420) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9420)))) severity failure;
    assert RAM(9421) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9421)))) severity failure;
    assert RAM(9422) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9422)))) severity failure;
    assert RAM(9423) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9423)))) severity failure;
    assert RAM(9424) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9424)))) severity failure;
    assert RAM(9425) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9425)))) severity failure;
    assert RAM(9426) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9426)))) severity failure;
    assert RAM(9427) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9427)))) severity failure;
    assert RAM(9428) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9428)))) severity failure;
    assert RAM(9429) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9429)))) severity failure;
    assert RAM(9430) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9430)))) severity failure;
    assert RAM(9431) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9431)))) severity failure;
    assert RAM(9432) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9432)))) severity failure;
    assert RAM(9433) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9433)))) severity failure;
    assert RAM(9434) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9434)))) severity failure;
    assert RAM(9435) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9435)))) severity failure;
    assert RAM(9436) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9436)))) severity failure;
    assert RAM(9437) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9437)))) severity failure;
    assert RAM(9438) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9438)))) severity failure;
    assert RAM(9439) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9439)))) severity failure;
    assert RAM(9440) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9440)))) severity failure;
    assert RAM(9441) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9441)))) severity failure;
    assert RAM(9442) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9442)))) severity failure;
    assert RAM(9443) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9443)))) severity failure;
    assert RAM(9444) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9444)))) severity failure;
    assert RAM(9445) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9445)))) severity failure;
    assert RAM(9446) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9446)))) severity failure;
    assert RAM(9447) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9447)))) severity failure;
    assert RAM(9448) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9448)))) severity failure;
    assert RAM(9449) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9449)))) severity failure;
    assert RAM(9450) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9450)))) severity failure;
    assert RAM(9451) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9451)))) severity failure;
    assert RAM(9452) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9452)))) severity failure;
    assert RAM(9453) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9453)))) severity failure;
    assert RAM(9454) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9454)))) severity failure;
    assert RAM(9455) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9455)))) severity failure;
    assert RAM(9456) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9456)))) severity failure;
    assert RAM(9457) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9457)))) severity failure;
    assert RAM(9458) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9458)))) severity failure;
    assert RAM(9459) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9459)))) severity failure;
    assert RAM(9460) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9460)))) severity failure;
    assert RAM(9461) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9461)))) severity failure;
    assert RAM(9462) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9462)))) severity failure;
    assert RAM(9463) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9463)))) severity failure;
    assert RAM(9464) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9464)))) severity failure;
    assert RAM(9465) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9465)))) severity failure;
    assert RAM(9466) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9466)))) severity failure;
    assert RAM(9467) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9467)))) severity failure;
    assert RAM(9468) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9468)))) severity failure;
    assert RAM(9469) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9469)))) severity failure;
    assert RAM(9470) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9470)))) severity failure;
    assert RAM(9471) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9471)))) severity failure;
    assert RAM(9472) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9472)))) severity failure;
    assert RAM(9473) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9473)))) severity failure;
    assert RAM(9474) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9474)))) severity failure;
    assert RAM(9475) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9475)))) severity failure;
    assert RAM(9476) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9476)))) severity failure;
    assert RAM(9477) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9477)))) severity failure;
    assert RAM(9478) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9478)))) severity failure;
    assert RAM(9479) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9479)))) severity failure;
    assert RAM(9480) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9480)))) severity failure;
    assert RAM(9481) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9481)))) severity failure;
    assert RAM(9482) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9482)))) severity failure;
    assert RAM(9483) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9483)))) severity failure;
    assert RAM(9484) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9484)))) severity failure;
    assert RAM(9485) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9485)))) severity failure;
    assert RAM(9486) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9486)))) severity failure;
    assert RAM(9487) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9487)))) severity failure;
    assert RAM(9488) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9488)))) severity failure;
    assert RAM(9489) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9489)))) severity failure;
    assert RAM(9490) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9490)))) severity failure;
    assert RAM(9491) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9491)))) severity failure;
    assert RAM(9492) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9492)))) severity failure;
    assert RAM(9493) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9493)))) severity failure;
    assert RAM(9494) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9494)))) severity failure;
    assert RAM(9495) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9495)))) severity failure;
    assert RAM(9496) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9496)))) severity failure;
    assert RAM(9497) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9497)))) severity failure;
    assert RAM(9498) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9498)))) severity failure;
    assert RAM(9499) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9499)))) severity failure;
    assert RAM(9500) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9500)))) severity failure;
    assert RAM(9501) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9501)))) severity failure;
    assert RAM(9502) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9502)))) severity failure;
    assert RAM(9503) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9503)))) severity failure;
    assert RAM(9504) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9504)))) severity failure;
    assert RAM(9505) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9505)))) severity failure;
    assert RAM(9506) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9506)))) severity failure;
    assert RAM(9507) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9507)))) severity failure;
    assert RAM(9508) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9508)))) severity failure;
    assert RAM(9509) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9509)))) severity failure;
    assert RAM(9510) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9510)))) severity failure;
    assert RAM(9511) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9511)))) severity failure;
    assert RAM(9512) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9512)))) severity failure;
    assert RAM(9513) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9513)))) severity failure;
    assert RAM(9514) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9514)))) severity failure;
    assert RAM(9515) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9515)))) severity failure;
    assert RAM(9516) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9516)))) severity failure;
    assert RAM(9517) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9517)))) severity failure;
    assert RAM(9518) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9518)))) severity failure;
    assert RAM(9519) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9519)))) severity failure;
    assert RAM(9520) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9520)))) severity failure;
    assert RAM(9521) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9521)))) severity failure;
    assert RAM(9522) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9522)))) severity failure;
    assert RAM(9523) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9523)))) severity failure;
    assert RAM(9524) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9524)))) severity failure;
    assert RAM(9525) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9525)))) severity failure;
    assert RAM(9526) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9526)))) severity failure;
    assert RAM(9527) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9527)))) severity failure;
    assert RAM(9528) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9528)))) severity failure;
    assert RAM(9529) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9529)))) severity failure;
    assert RAM(9530) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9530)))) severity failure;
    assert RAM(9531) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9531)))) severity failure;
    assert RAM(9532) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9532)))) severity failure;
    assert RAM(9533) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9533)))) severity failure;
    assert RAM(9534) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9534)))) severity failure;
    assert RAM(9535) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9535)))) severity failure;
    assert RAM(9536) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9536)))) severity failure;
    assert RAM(9537) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9537)))) severity failure;
    assert RAM(9538) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9538)))) severity failure;
    assert RAM(9539) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9539)))) severity failure;
    assert RAM(9540) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9540)))) severity failure;
    assert RAM(9541) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9541)))) severity failure;
    assert RAM(9542) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9542)))) severity failure;
    assert RAM(9543) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9543)))) severity failure;
    assert RAM(9544) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9544)))) severity failure;
    assert RAM(9545) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9545)))) severity failure;
    assert RAM(9546) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9546)))) severity failure;
    assert RAM(9547) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9547)))) severity failure;
    assert RAM(9548) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9548)))) severity failure;
    assert RAM(9549) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9549)))) severity failure;
    assert RAM(9550) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9550)))) severity failure;
    assert RAM(9551) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9551)))) severity failure;
    assert RAM(9552) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9552)))) severity failure;
    assert RAM(9553) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9553)))) severity failure;
    assert RAM(9554) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9554)))) severity failure;
    assert RAM(9555) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9555)))) severity failure;
    assert RAM(9556) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9556)))) severity failure;
    assert RAM(9557) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9557)))) severity failure;
    assert RAM(9558) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9558)))) severity failure;
    assert RAM(9559) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9559)))) severity failure;
    assert RAM(9560) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9560)))) severity failure;
    assert RAM(9561) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9561)))) severity failure;
    assert RAM(9562) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9562)))) severity failure;
    assert RAM(9563) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9563)))) severity failure;
    assert RAM(9564) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9564)))) severity failure;
    assert RAM(9565) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9565)))) severity failure;
    assert RAM(9566) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9566)))) severity failure;
    assert RAM(9567) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9567)))) severity failure;
    assert RAM(9568) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9568)))) severity failure;
    assert RAM(9569) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9569)))) severity failure;
    assert RAM(9570) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9570)))) severity failure;
    assert RAM(9571) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9571)))) severity failure;
    assert RAM(9572) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9572)))) severity failure;
    assert RAM(9573) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9573)))) severity failure;
    assert RAM(9574) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9574)))) severity failure;
    assert RAM(9575) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9575)))) severity failure;
    assert RAM(9576) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9576)))) severity failure;
    assert RAM(9577) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9577)))) severity failure;
    assert RAM(9578) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9578)))) severity failure;
    assert RAM(9579) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9579)))) severity failure;
    assert RAM(9580) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9580)))) severity failure;
    assert RAM(9581) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9581)))) severity failure;
    assert RAM(9582) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9582)))) severity failure;
    assert RAM(9583) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9583)))) severity failure;
    assert RAM(9584) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9584)))) severity failure;
    assert RAM(9585) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9585)))) severity failure;
    assert RAM(9586) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9586)))) severity failure;
    assert RAM(9587) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9587)))) severity failure;
    assert RAM(9588) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9588)))) severity failure;
    assert RAM(9589) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9589)))) severity failure;
    assert RAM(9590) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9590)))) severity failure;
    assert RAM(9591) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9591)))) severity failure;
    assert RAM(9592) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9592)))) severity failure;
    assert RAM(9593) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9593)))) severity failure;
    assert RAM(9594) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9594)))) severity failure;
    assert RAM(9595) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9595)))) severity failure;
    assert RAM(9596) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9596)))) severity failure;
    assert RAM(9597) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9597)))) severity failure;
    assert RAM(9598) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9598)))) severity failure;
    assert RAM(9599) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9599)))) severity failure;
    assert RAM(9600) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9600)))) severity failure;
    assert RAM(9601) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9601)))) severity failure;
    assert RAM(9602) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9602)))) severity failure;
    assert RAM(9603) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9603)))) severity failure;
    assert RAM(9604) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9604)))) severity failure;
    assert RAM(9605) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9605)))) severity failure;
    assert RAM(9606) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9606)))) severity failure;
    assert RAM(9607) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9607)))) severity failure;
    assert RAM(9608) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9608)))) severity failure;
    assert RAM(9609) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9609)))) severity failure;
    assert RAM(9610) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9610)))) severity failure;
    assert RAM(9611) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9611)))) severity failure;
    assert RAM(9612) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9612)))) severity failure;
    assert RAM(9613) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9613)))) severity failure;
    assert RAM(9614) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9614)))) severity failure;
    assert RAM(9615) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9615)))) severity failure;
    assert RAM(9616) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9616)))) severity failure;
    assert RAM(9617) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9617)))) severity failure;
    assert RAM(9618) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9618)))) severity failure;
    assert RAM(9619) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9619)))) severity failure;
    assert RAM(9620) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9620)))) severity failure;
    assert RAM(9621) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9621)))) severity failure;
    assert RAM(9622) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9622)))) severity failure;
    assert RAM(9623) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9623)))) severity failure;
    assert RAM(9624) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9624)))) severity failure;
    assert RAM(9625) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9625)))) severity failure;
    assert RAM(9626) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9626)))) severity failure;
    assert RAM(9627) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9627)))) severity failure;
    assert RAM(9628) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9628)))) severity failure;
    assert RAM(9629) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9629)))) severity failure;
    assert RAM(9630) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9630)))) severity failure;
    assert RAM(9631) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9631)))) severity failure;
    assert RAM(9632) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9632)))) severity failure;
    assert RAM(9633) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9633)))) severity failure;
    assert RAM(9634) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9634)))) severity failure;
    assert RAM(9635) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9635)))) severity failure;
    assert RAM(9636) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9636)))) severity failure;
    assert RAM(9637) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9637)))) severity failure;
    assert RAM(9638) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9638)))) severity failure;
    assert RAM(9639) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9639)))) severity failure;
    assert RAM(9640) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9640)))) severity failure;
    assert RAM(9641) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9641)))) severity failure;
    assert RAM(9642) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9642)))) severity failure;
    assert RAM(9643) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9643)))) severity failure;
    assert RAM(9644) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9644)))) severity failure;
    assert RAM(9645) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9645)))) severity failure;
    assert RAM(9646) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9646)))) severity failure;
    assert RAM(9647) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9647)))) severity failure;
    assert RAM(9648) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9648)))) severity failure;
    assert RAM(9649) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9649)))) severity failure;
    assert RAM(9650) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9650)))) severity failure;
    assert RAM(9651) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9651)))) severity failure;
    assert RAM(9652) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9652)))) severity failure;
    assert RAM(9653) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9653)))) severity failure;
    assert RAM(9654) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9654)))) severity failure;
    assert RAM(9655) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9655)))) severity failure;
    assert RAM(9656) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9656)))) severity failure;
    assert RAM(9657) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9657)))) severity failure;
    assert RAM(9658) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9658)))) severity failure;
    assert RAM(9659) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9659)))) severity failure;
    assert RAM(9660) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9660)))) severity failure;
    assert RAM(9661) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9661)))) severity failure;
    assert RAM(9662) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9662)))) severity failure;
    assert RAM(9663) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9663)))) severity failure;
    assert RAM(9664) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9664)))) severity failure;
    assert RAM(9665) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9665)))) severity failure;
    assert RAM(9666) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9666)))) severity failure;
    assert RAM(9667) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9667)))) severity failure;
    assert RAM(9668) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9668)))) severity failure;
    assert RAM(9669) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9669)))) severity failure;
    assert RAM(9670) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9670)))) severity failure;
    assert RAM(9671) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9671)))) severity failure;
    assert RAM(9672) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9672)))) severity failure;
    assert RAM(9673) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9673)))) severity failure;
    assert RAM(9674) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9674)))) severity failure;
    assert RAM(9675) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9675)))) severity failure;
    assert RAM(9676) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9676)))) severity failure;
    assert RAM(9677) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9677)))) severity failure;
    assert RAM(9678) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9678)))) severity failure;
    assert RAM(9679) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9679)))) severity failure;
    assert RAM(9680) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9680)))) severity failure;
    assert RAM(9681) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9681)))) severity failure;
    assert RAM(9682) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9682)))) severity failure;
    assert RAM(9683) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9683)))) severity failure;
    assert RAM(9684) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9684)))) severity failure;
    assert RAM(9685) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9685)))) severity failure;
    assert RAM(9686) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9686)))) severity failure;
    assert RAM(9687) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9687)))) severity failure;
    assert RAM(9688) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9688)))) severity failure;
    assert RAM(9689) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9689)))) severity failure;
    assert RAM(9690) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9690)))) severity failure;
    assert RAM(9691) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9691)))) severity failure;
    assert RAM(9692) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9692)))) severity failure;
    assert RAM(9693) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9693)))) severity failure;
    assert RAM(9694) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9694)))) severity failure;
    assert RAM(9695) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9695)))) severity failure;
    assert RAM(9696) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9696)))) severity failure;
    assert RAM(9697) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9697)))) severity failure;
    assert RAM(9698) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9698)))) severity failure;
    assert RAM(9699) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9699)))) severity failure;
    assert RAM(9700) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9700)))) severity failure;
    assert RAM(9701) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9701)))) severity failure;
    assert RAM(9702) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9702)))) severity failure;
    assert RAM(9703) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9703)))) severity failure;
    assert RAM(9704) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9704)))) severity failure;
    assert RAM(9705) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9705)))) severity failure;
    assert RAM(9706) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9706)))) severity failure;
    assert RAM(9707) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9707)))) severity failure;
    assert RAM(9708) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9708)))) severity failure;
    assert RAM(9709) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9709)))) severity failure;
    assert RAM(9710) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9710)))) severity failure;
    assert RAM(9711) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9711)))) severity failure;
    assert RAM(9712) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9712)))) severity failure;
    assert RAM(9713) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9713)))) severity failure;
    assert RAM(9714) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9714)))) severity failure;
    assert RAM(9715) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9715)))) severity failure;
    assert RAM(9716) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9716)))) severity failure;
    assert RAM(9717) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9717)))) severity failure;
    assert RAM(9718) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9718)))) severity failure;
    assert RAM(9719) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9719)))) severity failure;
    assert RAM(9720) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9720)))) severity failure;
    assert RAM(9721) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9721)))) severity failure;
    assert RAM(9722) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9722)))) severity failure;
    assert RAM(9723) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9723)))) severity failure;
    assert RAM(9724) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9724)))) severity failure;
    assert RAM(9725) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9725)))) severity failure;
    assert RAM(9726) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9726)))) severity failure;
    assert RAM(9727) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9727)))) severity failure;
    assert RAM(9728) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9728)))) severity failure;
    assert RAM(9729) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9729)))) severity failure;
    assert RAM(9730) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9730)))) severity failure;
    assert RAM(9731) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9731)))) severity failure;
    assert RAM(9732) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9732)))) severity failure;
    assert RAM(9733) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9733)))) severity failure;
    assert RAM(9734) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9734)))) severity failure;
    assert RAM(9735) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9735)))) severity failure;
    assert RAM(9736) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9736)))) severity failure;
    assert RAM(9737) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9737)))) severity failure;
    assert RAM(9738) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9738)))) severity failure;
    assert RAM(9739) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9739)))) severity failure;
    assert RAM(9740) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9740)))) severity failure;
    assert RAM(9741) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9741)))) severity failure;
    assert RAM(9742) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9742)))) severity failure;
    assert RAM(9743) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9743)))) severity failure;
    assert RAM(9744) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9744)))) severity failure;
    assert RAM(9745) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9745)))) severity failure;
    assert RAM(9746) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9746)))) severity failure;
    assert RAM(9747) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9747)))) severity failure;
    assert RAM(9748) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9748)))) severity failure;
    assert RAM(9749) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9749)))) severity failure;
    assert RAM(9750) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9750)))) severity failure;
    assert RAM(9751) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9751)))) severity failure;
    assert RAM(9752) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9752)))) severity failure;
    assert RAM(9753) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9753)))) severity failure;
    assert RAM(9754) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9754)))) severity failure;
    assert RAM(9755) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9755)))) severity failure;
    assert RAM(9756) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9756)))) severity failure;
    assert RAM(9757) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9757)))) severity failure;
    assert RAM(9758) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9758)))) severity failure;
    assert RAM(9759) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9759)))) severity failure;
    assert RAM(9760) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9760)))) severity failure;
    assert RAM(9761) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9761)))) severity failure;
    assert RAM(9762) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9762)))) severity failure;
    assert RAM(9763) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9763)))) severity failure;
    assert RAM(9764) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9764)))) severity failure;
    assert RAM(9765) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9765)))) severity failure;
    assert RAM(9766) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9766)))) severity failure;
    assert RAM(9767) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9767)))) severity failure;
    assert RAM(9768) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9768)))) severity failure;
    assert RAM(9769) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9769)))) severity failure;
    assert RAM(9770) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9770)))) severity failure;
    assert RAM(9771) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9771)))) severity failure;
    assert RAM(9772) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9772)))) severity failure;
    assert RAM(9773) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9773)))) severity failure;
    assert RAM(9774) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9774)))) severity failure;
    assert RAM(9775) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9775)))) severity failure;
    assert RAM(9776) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9776)))) severity failure;
    assert RAM(9777) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9777)))) severity failure;
    assert RAM(9778) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9778)))) severity failure;
    assert RAM(9779) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9779)))) severity failure;
    assert RAM(9780) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9780)))) severity failure;
    assert RAM(9781) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9781)))) severity failure;
    assert RAM(9782) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9782)))) severity failure;
    assert RAM(9783) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9783)))) severity failure;
    assert RAM(9784) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9784)))) severity failure;
    assert RAM(9785) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9785)))) severity failure;
    assert RAM(9786) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9786)))) severity failure;
    assert RAM(9787) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9787)))) severity failure;
    assert RAM(9788) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9788)))) severity failure;
    assert RAM(9789) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9789)))) severity failure;
    assert RAM(9790) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9790)))) severity failure;
    assert RAM(9791) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9791)))) severity failure;
    assert RAM(9792) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9792)))) severity failure;
    assert RAM(9793) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9793)))) severity failure;
    assert RAM(9794) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9794)))) severity failure;
    assert RAM(9795) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9795)))) severity failure;
    assert RAM(9796) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9796)))) severity failure;
    assert RAM(9797) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9797)))) severity failure;
    assert RAM(9798) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9798)))) severity failure;
    assert RAM(9799) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9799)))) severity failure;
    assert RAM(9800) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9800)))) severity failure;
    assert RAM(9801) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9801)))) severity failure;
    assert RAM(9802) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9802)))) severity failure;
    assert RAM(9803) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9803)))) severity failure;
    assert RAM(9804) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9804)))) severity failure;
    assert RAM(9805) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9805)))) severity failure;
    assert RAM(9806) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9806)))) severity failure;
    assert RAM(9807) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9807)))) severity failure;
    assert RAM(9808) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9808)))) severity failure;
    assert RAM(9809) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9809)))) severity failure;
    assert RAM(9810) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9810)))) severity failure;
    assert RAM(9811) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9811)))) severity failure;
    assert RAM(9812) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9812)))) severity failure;
    assert RAM(9813) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9813)))) severity failure;
    assert RAM(9814) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9814)))) severity failure;
    assert RAM(9815) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9815)))) severity failure;
    assert RAM(9816) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9816)))) severity failure;
    assert RAM(9817) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9817)))) severity failure;
    assert RAM(9818) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9818)))) severity failure;
    assert RAM(9819) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9819)))) severity failure;
    assert RAM(9820) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9820)))) severity failure;
    assert RAM(9821) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9821)))) severity failure;
    assert RAM(9822) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9822)))) severity failure;
    assert RAM(9823) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9823)))) severity failure;
    assert RAM(9824) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9824)))) severity failure;
    assert RAM(9825) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9825)))) severity failure;
    assert RAM(9826) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9826)))) severity failure;
    assert RAM(9827) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9827)))) severity failure;
    assert RAM(9828) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9828)))) severity failure;
    assert RAM(9829) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9829)))) severity failure;
    assert RAM(9830) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9830)))) severity failure;
    assert RAM(9831) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9831)))) severity failure;
    assert RAM(9832) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9832)))) severity failure;
    assert RAM(9833) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9833)))) severity failure;
    assert RAM(9834) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9834)))) severity failure;
    assert RAM(9835) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9835)))) severity failure;
    assert RAM(9836) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9836)))) severity failure;
    assert RAM(9837) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9837)))) severity failure;
    assert RAM(9838) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9838)))) severity failure;
    assert RAM(9839) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9839)))) severity failure;
    assert RAM(9840) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9840)))) severity failure;
    assert RAM(9841) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9841)))) severity failure;
    assert RAM(9842) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9842)))) severity failure;
    assert RAM(9843) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9843)))) severity failure;
    assert RAM(9844) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9844)))) severity failure;
    assert RAM(9845) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9845)))) severity failure;
    assert RAM(9846) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9846)))) severity failure;
    assert RAM(9847) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9847)))) severity failure;
    assert RAM(9848) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9848)))) severity failure;
    assert RAM(9849) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9849)))) severity failure;
    assert RAM(9850) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9850)))) severity failure;
    assert RAM(9851) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9851)))) severity failure;
    assert RAM(9852) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9852)))) severity failure;
    assert RAM(9853) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9853)))) severity failure;
    assert RAM(9854) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9854)))) severity failure;
    assert RAM(9855) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9855)))) severity failure;
    assert RAM(9856) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9856)))) severity failure;
    assert RAM(9857) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9857)))) severity failure;
    assert RAM(9858) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9858)))) severity failure;
    assert RAM(9859) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9859)))) severity failure;
    assert RAM(9860) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9860)))) severity failure;
    assert RAM(9861) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9861)))) severity failure;
    assert RAM(9862) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9862)))) severity failure;
    assert RAM(9863) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9863)))) severity failure;
    assert RAM(9864) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9864)))) severity failure;
    assert RAM(9865) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9865)))) severity failure;
    assert RAM(9866) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9866)))) severity failure;
    assert RAM(9867) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9867)))) severity failure;
    assert RAM(9868) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9868)))) severity failure;
    assert RAM(9869) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9869)))) severity failure;
    assert RAM(9870) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9870)))) severity failure;
    assert RAM(9871) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9871)))) severity failure;
    assert RAM(9872) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9872)))) severity failure;
    assert RAM(9873) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9873)))) severity failure;
    assert RAM(9874) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9874)))) severity failure;
    assert RAM(9875) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9875)))) severity failure;
    assert RAM(9876) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9876)))) severity failure;
    assert RAM(9877) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9877)))) severity failure;
    assert RAM(9878) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9878)))) severity failure;
    assert RAM(9879) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9879)))) severity failure;
    assert RAM(9880) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9880)))) severity failure;
    assert RAM(9881) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9881)))) severity failure;
    assert RAM(9882) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9882)))) severity failure;
    assert RAM(9883) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9883)))) severity failure;
    assert RAM(9884) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9884)))) severity failure;
    assert RAM(9885) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9885)))) severity failure;
    assert RAM(9886) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9886)))) severity failure;
    assert RAM(9887) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9887)))) severity failure;
    assert RAM(9888) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9888)))) severity failure;
    assert RAM(9889) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9889)))) severity failure;
    assert RAM(9890) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9890)))) severity failure;
    assert RAM(9891) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9891)))) severity failure;
    assert RAM(9892) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9892)))) severity failure;
    assert RAM(9893) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9893)))) severity failure;
    assert RAM(9894) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9894)))) severity failure;
    assert RAM(9895) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9895)))) severity failure;
    assert RAM(9896) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9896)))) severity failure;
    assert RAM(9897) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9897)))) severity failure;
    assert RAM(9898) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9898)))) severity failure;
    assert RAM(9899) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9899)))) severity failure;
    assert RAM(9900) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9900)))) severity failure;
    assert RAM(9901) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9901)))) severity failure;
    assert RAM(9902) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9902)))) severity failure;
    assert RAM(9903) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9903)))) severity failure;
    assert RAM(9904) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9904)))) severity failure;
    assert RAM(9905) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9905)))) severity failure;
    assert RAM(9906) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9906)))) severity failure;
    assert RAM(9907) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9907)))) severity failure;
    assert RAM(9908) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9908)))) severity failure;
    assert RAM(9909) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9909)))) severity failure;
    assert RAM(9910) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9910)))) severity failure;
    assert RAM(9911) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9911)))) severity failure;
    assert RAM(9912) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9912)))) severity failure;
    assert RAM(9913) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9913)))) severity failure;
    assert RAM(9914) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9914)))) severity failure;
    assert RAM(9915) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9915)))) severity failure;
    assert RAM(9916) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9916)))) severity failure;
    assert RAM(9917) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9917)))) severity failure;
    assert RAM(9918) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9918)))) severity failure;
    assert RAM(9919) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9919)))) severity failure;
    assert RAM(9920) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9920)))) severity failure;
    assert RAM(9921) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9921)))) severity failure;
    assert RAM(9922) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9922)))) severity failure;
    assert RAM(9923) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9923)))) severity failure;
    assert RAM(9924) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9924)))) severity failure;
    assert RAM(9925) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9925)))) severity failure;
    assert RAM(9926) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9926)))) severity failure;
    assert RAM(9927) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9927)))) severity failure;
    assert RAM(9928) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9928)))) severity failure;
    assert RAM(9929) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9929)))) severity failure;
    assert RAM(9930) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9930)))) severity failure;
    assert RAM(9931) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9931)))) severity failure;
    assert RAM(9932) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9932)))) severity failure;
    assert RAM(9933) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9933)))) severity failure;
    assert RAM(9934) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9934)))) severity failure;
    assert RAM(9935) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9935)))) severity failure;
    assert RAM(9936) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9936)))) severity failure;
    assert RAM(9937) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9937)))) severity failure;
    assert RAM(9938) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9938)))) severity failure;
    assert RAM(9939) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9939)))) severity failure;
    assert RAM(9940) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9940)))) severity failure;
    assert RAM(9941) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9941)))) severity failure;
    assert RAM(9942) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9942)))) severity failure;
    assert RAM(9943) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9943)))) severity failure;
    assert RAM(9944) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9944)))) severity failure;
    assert RAM(9945) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9945)))) severity failure;
    assert RAM(9946) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9946)))) severity failure;
    assert RAM(9947) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9947)))) severity failure;
    assert RAM(9948) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9948)))) severity failure;
    assert RAM(9949) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9949)))) severity failure;
    assert RAM(9950) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9950)))) severity failure;
    assert RAM(9951) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9951)))) severity failure;
    assert RAM(9952) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9952)))) severity failure;
    assert RAM(9953) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9953)))) severity failure;
    assert RAM(9954) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9954)))) severity failure;
    assert RAM(9955) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9955)))) severity failure;
    assert RAM(9956) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9956)))) severity failure;
    assert RAM(9957) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9957)))) severity failure;
    assert RAM(9958) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9958)))) severity failure;
    assert RAM(9959) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9959)))) severity failure;
    assert RAM(9960) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9960)))) severity failure;
    assert RAM(9961) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9961)))) severity failure;
    assert RAM(9962) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9962)))) severity failure;
    assert RAM(9963) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9963)))) severity failure;
    assert RAM(9964) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9964)))) severity failure;
    assert RAM(9965) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9965)))) severity failure;
    assert RAM(9966) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9966)))) severity failure;
    assert RAM(9967) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9967)))) severity failure;
    assert RAM(9968) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9968)))) severity failure;
    assert RAM(9969) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9969)))) severity failure;
    assert RAM(9970) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9970)))) severity failure;
    assert RAM(9971) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9971)))) severity failure;
    assert RAM(9972) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9972)))) severity failure;
    assert RAM(9973) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9973)))) severity failure;
    assert RAM(9974) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9974)))) severity failure;
    assert RAM(9975) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9975)))) severity failure;
    assert RAM(9976) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9976)))) severity failure;
    assert RAM(9977) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9977)))) severity failure;
    assert RAM(9978) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9978)))) severity failure;
    assert RAM(9979) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9979)))) severity failure;
    assert RAM(9980) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9980)))) severity failure;
    assert RAM(9981) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9981)))) severity failure;
    assert RAM(9982) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9982)))) severity failure;
    assert RAM(9983) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9983)))) severity failure;
    assert RAM(9984) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9984)))) severity failure;
    assert RAM(9985) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9985)))) severity failure;
    assert RAM(9986) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9986)))) severity failure;
    assert RAM(9987) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9987)))) severity failure;
    assert RAM(9988) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9988)))) severity failure;
    assert RAM(9989) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9989)))) severity failure;
    assert RAM(9990) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9990)))) severity failure;
    assert RAM(9991) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9991)))) severity failure;
    assert RAM(9992) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9992)))) severity failure;
    assert RAM(9993) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9993)))) severity failure;
    assert RAM(9994) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9994)))) severity failure;
    assert RAM(9995) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9995)))) severity failure;
    assert RAM(9996) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9996)))) severity failure;
    assert RAM(9997) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9997)))) severity failure;
    assert RAM(9998) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(9998)))) severity failure;
    assert RAM(9999) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(9999)))) severity failure;
    assert RAM(10000) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10000)))) severity failure;
    assert RAM(10001) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10001)))) severity failure;
    assert RAM(10002) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10002)))) severity failure;
    assert RAM(10003) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10003)))) severity failure;
    assert RAM(10004) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10004)))) severity failure;
    assert RAM(10005) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10005)))) severity failure;
    assert RAM(10006) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10006)))) severity failure;
    assert RAM(10007) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10007)))) severity failure;
    assert RAM(10008) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10008)))) severity failure;
    assert RAM(10009) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10009)))) severity failure;
    assert RAM(10010) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10010)))) severity failure;
    assert RAM(10011) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10011)))) severity failure;
    assert RAM(10012) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10012)))) severity failure;
    assert RAM(10013) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10013)))) severity failure;
    assert RAM(10014) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10014)))) severity failure;
    assert RAM(10015) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10015)))) severity failure;
    assert RAM(10016) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10016)))) severity failure;
    assert RAM(10017) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10017)))) severity failure;
    assert RAM(10018) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10018)))) severity failure;
    assert RAM(10019) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10019)))) severity failure;
    assert RAM(10020) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10020)))) severity failure;
    assert RAM(10021) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10021)))) severity failure;
    assert RAM(10022) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10022)))) severity failure;
    assert RAM(10023) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10023)))) severity failure;
    assert RAM(10024) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10024)))) severity failure;
    assert RAM(10025) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10025)))) severity failure;
    assert RAM(10026) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10026)))) severity failure;
    assert RAM(10027) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10027)))) severity failure;
    assert RAM(10028) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10028)))) severity failure;
    assert RAM(10029) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10029)))) severity failure;
    assert RAM(10030) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10030)))) severity failure;
    assert RAM(10031) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10031)))) severity failure;
    assert RAM(10032) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10032)))) severity failure;
    assert RAM(10033) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10033)))) severity failure;
    assert RAM(10034) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10034)))) severity failure;
    assert RAM(10035) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10035)))) severity failure;
    assert RAM(10036) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10036)))) severity failure;
    assert RAM(10037) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10037)))) severity failure;
    assert RAM(10038) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10038)))) severity failure;
    assert RAM(10039) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10039)))) severity failure;
    assert RAM(10040) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10040)))) severity failure;
    assert RAM(10041) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10041)))) severity failure;
    assert RAM(10042) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10042)))) severity failure;
    assert RAM(10043) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10043)))) severity failure;
    assert RAM(10044) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10044)))) severity failure;
    assert RAM(10045) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10045)))) severity failure;
    assert RAM(10046) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10046)))) severity failure;
    assert RAM(10047) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10047)))) severity failure;
    assert RAM(10048) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10048)))) severity failure;
    assert RAM(10049) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10049)))) severity failure;
    assert RAM(10050) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10050)))) severity failure;
    assert RAM(10051) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10051)))) severity failure;
    assert RAM(10052) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10052)))) severity failure;
    assert RAM(10053) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10053)))) severity failure;
    assert RAM(10054) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10054)))) severity failure;
    assert RAM(10055) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10055)))) severity failure;
    assert RAM(10056) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10056)))) severity failure;
    assert RAM(10057) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10057)))) severity failure;
    assert RAM(10058) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10058)))) severity failure;
    assert RAM(10059) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10059)))) severity failure;
    assert RAM(10060) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10060)))) severity failure;
    assert RAM(10061) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10061)))) severity failure;
    assert RAM(10062) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10062)))) severity failure;
    assert RAM(10063) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10063)))) severity failure;
    assert RAM(10064) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10064)))) severity failure;
    assert RAM(10065) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10065)))) severity failure;
    assert RAM(10066) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10066)))) severity failure;
    assert RAM(10067) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10067)))) severity failure;
    assert RAM(10068) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10068)))) severity failure;
    assert RAM(10069) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10069)))) severity failure;
    assert RAM(10070) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10070)))) severity failure;
    assert RAM(10071) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10071)))) severity failure;
    assert RAM(10072) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10072)))) severity failure;
    assert RAM(10073) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10073)))) severity failure;
    assert RAM(10074) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10074)))) severity failure;
    assert RAM(10075) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10075)))) severity failure;
    assert RAM(10076) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10076)))) severity failure;
    assert RAM(10077) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10077)))) severity failure;
    assert RAM(10078) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10078)))) severity failure;
    assert RAM(10079) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10079)))) severity failure;
    assert RAM(10080) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10080)))) severity failure;
    assert RAM(10081) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10081)))) severity failure;
    assert RAM(10082) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10082)))) severity failure;
    assert RAM(10083) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10083)))) severity failure;
    assert RAM(10084) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10084)))) severity failure;
    assert RAM(10085) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10085)))) severity failure;
    assert RAM(10086) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10086)))) severity failure;
    assert RAM(10087) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10087)))) severity failure;
    assert RAM(10088) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10088)))) severity failure;
    assert RAM(10089) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10089)))) severity failure;
    assert RAM(10090) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10090)))) severity failure;
    assert RAM(10091) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10091)))) severity failure;
    assert RAM(10092) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10092)))) severity failure;
    assert RAM(10093) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10093)))) severity failure;
    assert RAM(10094) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10094)))) severity failure;
    assert RAM(10095) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10095)))) severity failure;
    assert RAM(10096) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10096)))) severity failure;
    assert RAM(10097) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10097)))) severity failure;
    assert RAM(10098) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10098)))) severity failure;
    assert RAM(10099) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10099)))) severity failure;
    assert RAM(10100) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10100)))) severity failure;
    assert RAM(10101) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10101)))) severity failure;
    assert RAM(10102) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10102)))) severity failure;
    assert RAM(10103) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10103)))) severity failure;
    assert RAM(10104) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10104)))) severity failure;
    assert RAM(10105) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10105)))) severity failure;
    assert RAM(10106) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10106)))) severity failure;
    assert RAM(10107) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10107)))) severity failure;
    assert RAM(10108) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10108)))) severity failure;
    assert RAM(10109) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10109)))) severity failure;
    assert RAM(10110) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10110)))) severity failure;
    assert RAM(10111) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10111)))) severity failure;
    assert RAM(10112) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10112)))) severity failure;
    assert RAM(10113) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10113)))) severity failure;
    assert RAM(10114) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10114)))) severity failure;
    assert RAM(10115) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10115)))) severity failure;
    assert RAM(10116) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10116)))) severity failure;
    assert RAM(10117) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10117)))) severity failure;
    assert RAM(10118) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10118)))) severity failure;
    assert RAM(10119) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10119)))) severity failure;
    assert RAM(10120) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10120)))) severity failure;
    assert RAM(10121) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10121)))) severity failure;
    assert RAM(10122) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10122)))) severity failure;
    assert RAM(10123) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10123)))) severity failure;
    assert RAM(10124) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10124)))) severity failure;
    assert RAM(10125) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10125)))) severity failure;
    assert RAM(10126) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10126)))) severity failure;
    assert RAM(10127) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10127)))) severity failure;
    assert RAM(10128) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10128)))) severity failure;
    assert RAM(10129) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10129)))) severity failure;
    assert RAM(10130) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10130)))) severity failure;
    assert RAM(10131) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10131)))) severity failure;
    assert RAM(10132) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10132)))) severity failure;
    assert RAM(10133) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10133)))) severity failure;
    assert RAM(10134) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10134)))) severity failure;
    assert RAM(10135) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10135)))) severity failure;
    assert RAM(10136) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10136)))) severity failure;
    assert RAM(10137) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10137)))) severity failure;
    assert RAM(10138) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10138)))) severity failure;
    assert RAM(10139) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10139)))) severity failure;
    assert RAM(10140) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10140)))) severity failure;
    assert RAM(10141) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10141)))) severity failure;
    assert RAM(10142) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10142)))) severity failure;
    assert RAM(10143) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10143)))) severity failure;
    assert RAM(10144) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10144)))) severity failure;
    assert RAM(10145) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10145)))) severity failure;
    assert RAM(10146) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10146)))) severity failure;
    assert RAM(10147) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10147)))) severity failure;
    assert RAM(10148) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10148)))) severity failure;
    assert RAM(10149) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10149)))) severity failure;
    assert RAM(10150) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10150)))) severity failure;
    assert RAM(10151) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10151)))) severity failure;
    assert RAM(10152) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10152)))) severity failure;
    assert RAM(10153) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10153)))) severity failure;
    assert RAM(10154) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10154)))) severity failure;
    assert RAM(10155) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10155)))) severity failure;
    assert RAM(10156) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10156)))) severity failure;
    assert RAM(10157) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10157)))) severity failure;
    assert RAM(10158) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10158)))) severity failure;
    assert RAM(10159) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10159)))) severity failure;
    assert RAM(10160) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10160)))) severity failure;
    assert RAM(10161) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10161)))) severity failure;
    assert RAM(10162) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10162)))) severity failure;
    assert RAM(10163) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10163)))) severity failure;
    assert RAM(10164) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10164)))) severity failure;
    assert RAM(10165) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10165)))) severity failure;
    assert RAM(10166) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10166)))) severity failure;
    assert RAM(10167) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10167)))) severity failure;
    assert RAM(10168) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10168)))) severity failure;
    assert RAM(10169) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10169)))) severity failure;
    assert RAM(10170) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10170)))) severity failure;
    assert RAM(10171) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10171)))) severity failure;
    assert RAM(10172) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10172)))) severity failure;
    assert RAM(10173) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10173)))) severity failure;
    assert RAM(10174) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10174)))) severity failure;
    assert RAM(10175) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10175)))) severity failure;
    assert RAM(10176) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10176)))) severity failure;
    assert RAM(10177) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10177)))) severity failure;
    assert RAM(10178) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10178)))) severity failure;
    assert RAM(10179) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10179)))) severity failure;
    assert RAM(10180) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10180)))) severity failure;
    assert RAM(10181) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10181)))) severity failure;
    assert RAM(10182) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10182)))) severity failure;
    assert RAM(10183) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10183)))) severity failure;
    assert RAM(10184) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10184)))) severity failure;
    assert RAM(10185) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10185)))) severity failure;
    assert RAM(10186) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10186)))) severity failure;
    assert RAM(10187) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10187)))) severity failure;
    assert RAM(10188) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10188)))) severity failure;
    assert RAM(10189) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10189)))) severity failure;
    assert RAM(10190) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10190)))) severity failure;
    assert RAM(10191) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10191)))) severity failure;
    assert RAM(10192) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10192)))) severity failure;
    assert RAM(10193) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10193)))) severity failure;
    assert RAM(10194) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10194)))) severity failure;
    assert RAM(10195) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10195)))) severity failure;
    assert RAM(10196) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10196)))) severity failure;
    assert RAM(10197) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10197)))) severity failure;
    assert RAM(10198) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10198)))) severity failure;
    assert RAM(10199) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10199)))) severity failure;
    assert RAM(10200) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10200)))) severity failure;
    assert RAM(10201) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10201)))) severity failure;
    assert RAM(10202) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10202)))) severity failure;
    assert RAM(10203) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10203)))) severity failure;
    assert RAM(10204) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10204)))) severity failure;
    assert RAM(10205) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10205)))) severity failure;
    assert RAM(10206) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10206)))) severity failure;
    assert RAM(10207) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10207)))) severity failure;
    assert RAM(10208) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10208)))) severity failure;
    assert RAM(10209) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10209)))) severity failure;
    assert RAM(10210) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10210)))) severity failure;
    assert RAM(10211) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10211)))) severity failure;
    assert RAM(10212) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10212)))) severity failure;
    assert RAM(10213) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10213)))) severity failure;
    assert RAM(10214) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10214)))) severity failure;
    assert RAM(10215) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10215)))) severity failure;
    assert RAM(10216) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10216)))) severity failure;
    assert RAM(10217) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10217)))) severity failure;
    assert RAM(10218) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10218)))) severity failure;
    assert RAM(10219) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10219)))) severity failure;
    assert RAM(10220) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10220)))) severity failure;
    assert RAM(10221) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10221)))) severity failure;
    assert RAM(10222) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10222)))) severity failure;
    assert RAM(10223) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10223)))) severity failure;
    assert RAM(10224) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10224)))) severity failure;
    assert RAM(10225) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10225)))) severity failure;
    assert RAM(10226) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10226)))) severity failure;
    assert RAM(10227) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10227)))) severity failure;
    assert RAM(10228) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10228)))) severity failure;
    assert RAM(10229) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10229)))) severity failure;
    assert RAM(10230) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10230)))) severity failure;
    assert RAM(10231) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10231)))) severity failure;
    assert RAM(10232) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10232)))) severity failure;
    assert RAM(10233) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10233)))) severity failure;
    assert RAM(10234) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10234)))) severity failure;
    assert RAM(10235) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10235)))) severity failure;
    assert RAM(10236) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10236)))) severity failure;
    assert RAM(10237) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10237)))) severity failure;
    assert RAM(10238) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10238)))) severity failure;
    assert RAM(10239) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10239)))) severity failure;
    assert RAM(10240) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10240)))) severity failure;
    assert RAM(10241) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10241)))) severity failure;
    assert RAM(10242) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10242)))) severity failure;
    assert RAM(10243) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10243)))) severity failure;
    assert RAM(10244) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10244)))) severity failure;
    assert RAM(10245) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10245)))) severity failure;
    assert RAM(10246) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10246)))) severity failure;
    assert RAM(10247) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10247)))) severity failure;
    assert RAM(10248) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10248)))) severity failure;
    assert RAM(10249) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10249)))) severity failure;
    assert RAM(10250) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10250)))) severity failure;
    assert RAM(10251) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10251)))) severity failure;
    assert RAM(10252) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10252)))) severity failure;
    assert RAM(10253) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10253)))) severity failure;
    assert RAM(10254) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10254)))) severity failure;
    assert RAM(10255) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10255)))) severity failure;
    assert RAM(10256) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10256)))) severity failure;
    assert RAM(10257) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10257)))) severity failure;
    assert RAM(10258) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10258)))) severity failure;
    assert RAM(10259) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10259)))) severity failure;
    assert RAM(10260) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10260)))) severity failure;
    assert RAM(10261) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10261)))) severity failure;
    assert RAM(10262) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10262)))) severity failure;
    assert RAM(10263) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10263)))) severity failure;
    assert RAM(10264) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10264)))) severity failure;
    assert RAM(10265) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10265)))) severity failure;
    assert RAM(10266) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10266)))) severity failure;
    assert RAM(10267) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10267)))) severity failure;
    assert RAM(10268) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10268)))) severity failure;
    assert RAM(10269) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10269)))) severity failure;
    assert RAM(10270) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10270)))) severity failure;
    assert RAM(10271) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10271)))) severity failure;
    assert RAM(10272) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10272)))) severity failure;
    assert RAM(10273) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10273)))) severity failure;
    assert RAM(10274) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10274)))) severity failure;
    assert RAM(10275) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10275)))) severity failure;
    assert RAM(10276) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10276)))) severity failure;
    assert RAM(10277) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10277)))) severity failure;
    assert RAM(10278) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10278)))) severity failure;
    assert RAM(10279) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10279)))) severity failure;
    assert RAM(10280) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10280)))) severity failure;
    assert RAM(10281) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10281)))) severity failure;
    assert RAM(10282) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10282)))) severity failure;
    assert RAM(10283) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10283)))) severity failure;
    assert RAM(10284) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10284)))) severity failure;
    assert RAM(10285) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10285)))) severity failure;
    assert RAM(10286) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10286)))) severity failure;
    assert RAM(10287) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10287)))) severity failure;
    assert RAM(10288) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10288)))) severity failure;
    assert RAM(10289) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10289)))) severity failure;
    assert RAM(10290) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10290)))) severity failure;
    assert RAM(10291) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10291)))) severity failure;
    assert RAM(10292) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10292)))) severity failure;
    assert RAM(10293) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10293)))) severity failure;
    assert RAM(10294) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10294)))) severity failure;
    assert RAM(10295) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10295)))) severity failure;
    assert RAM(10296) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10296)))) severity failure;
    assert RAM(10297) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10297)))) severity failure;
    assert RAM(10298) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10298)))) severity failure;
    assert RAM(10299) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10299)))) severity failure;
    assert RAM(10300) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10300)))) severity failure;
    assert RAM(10301) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10301)))) severity failure;
    assert RAM(10302) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10302)))) severity failure;
    assert RAM(10303) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10303)))) severity failure;
    assert RAM(10304) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10304)))) severity failure;
    assert RAM(10305) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10305)))) severity failure;
    assert RAM(10306) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10306)))) severity failure;
    assert RAM(10307) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10307)))) severity failure;
    assert RAM(10308) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10308)))) severity failure;
    assert RAM(10309) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10309)))) severity failure;
    assert RAM(10310) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10310)))) severity failure;
    assert RAM(10311) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10311)))) severity failure;
    assert RAM(10312) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10312)))) severity failure;
    assert RAM(10313) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10313)))) severity failure;
    assert RAM(10314) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10314)))) severity failure;
    assert RAM(10315) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10315)))) severity failure;
    assert RAM(10316) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10316)))) severity failure;
    assert RAM(10317) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10317)))) severity failure;
    assert RAM(10318) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10318)))) severity failure;
    assert RAM(10319) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10319)))) severity failure;
    assert RAM(10320) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10320)))) severity failure;
    assert RAM(10321) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10321)))) severity failure;
    assert RAM(10322) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10322)))) severity failure;
    assert RAM(10323) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10323)))) severity failure;
    assert RAM(10324) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10324)))) severity failure;
    assert RAM(10325) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10325)))) severity failure;
    assert RAM(10326) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10326)))) severity failure;
    assert RAM(10327) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10327)))) severity failure;
    assert RAM(10328) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10328)))) severity failure;
    assert RAM(10329) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10329)))) severity failure;
    assert RAM(10330) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10330)))) severity failure;
    assert RAM(10331) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10331)))) severity failure;
    assert RAM(10332) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10332)))) severity failure;
    assert RAM(10333) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10333)))) severity failure;
    assert RAM(10334) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10334)))) severity failure;
    assert RAM(10335) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10335)))) severity failure;
    assert RAM(10336) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10336)))) severity failure;
    assert RAM(10337) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10337)))) severity failure;
    assert RAM(10338) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10338)))) severity failure;
    assert RAM(10339) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10339)))) severity failure;
    assert RAM(10340) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10340)))) severity failure;
    assert RAM(10341) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10341)))) severity failure;
    assert RAM(10342) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10342)))) severity failure;
    assert RAM(10343) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10343)))) severity failure;
    assert RAM(10344) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10344)))) severity failure;
    assert RAM(10345) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10345)))) severity failure;
    assert RAM(10346) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10346)))) severity failure;
    assert RAM(10347) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10347)))) severity failure;
    assert RAM(10348) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10348)))) severity failure;
    assert RAM(10349) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10349)))) severity failure;
    assert RAM(10350) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10350)))) severity failure;
    assert RAM(10351) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10351)))) severity failure;
    assert RAM(10352) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10352)))) severity failure;
    assert RAM(10353) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10353)))) severity failure;
    assert RAM(10354) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10354)))) severity failure;
    assert RAM(10355) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10355)))) severity failure;
    assert RAM(10356) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10356)))) severity failure;
    assert RAM(10357) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10357)))) severity failure;
    assert RAM(10358) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10358)))) severity failure;
    assert RAM(10359) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10359)))) severity failure;
    assert RAM(10360) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10360)))) severity failure;
    assert RAM(10361) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10361)))) severity failure;
    assert RAM(10362) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10362)))) severity failure;
    assert RAM(10363) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10363)))) severity failure;
    assert RAM(10364) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10364)))) severity failure;
    assert RAM(10365) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10365)))) severity failure;
    assert RAM(10366) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10366)))) severity failure;
    assert RAM(10367) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10367)))) severity failure;
    assert RAM(10368) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10368)))) severity failure;
    assert RAM(10369) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10369)))) severity failure;
    assert RAM(10370) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10370)))) severity failure;
    assert RAM(10371) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10371)))) severity failure;
    assert RAM(10372) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10372)))) severity failure;
    assert RAM(10373) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10373)))) severity failure;
    assert RAM(10374) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10374)))) severity failure;
    assert RAM(10375) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10375)))) severity failure;
    assert RAM(10376) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10376)))) severity failure;
    assert RAM(10377) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10377)))) severity failure;
    assert RAM(10378) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10378)))) severity failure;
    assert RAM(10379) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10379)))) severity failure;
    assert RAM(10380) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10380)))) severity failure;
    assert RAM(10381) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10381)))) severity failure;
    assert RAM(10382) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10382)))) severity failure;
    assert RAM(10383) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10383)))) severity failure;
    assert RAM(10384) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10384)))) severity failure;
    assert RAM(10385) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10385)))) severity failure;
    assert RAM(10386) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10386)))) severity failure;
    assert RAM(10387) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10387)))) severity failure;
    assert RAM(10388) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10388)))) severity failure;
    assert RAM(10389) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10389)))) severity failure;
    assert RAM(10390) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10390)))) severity failure;
    assert RAM(10391) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10391)))) severity failure;
    assert RAM(10392) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10392)))) severity failure;
    assert RAM(10393) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10393)))) severity failure;
    assert RAM(10394) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10394)))) severity failure;
    assert RAM(10395) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10395)))) severity failure;
    assert RAM(10396) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10396)))) severity failure;
    assert RAM(10397) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10397)))) severity failure;
    assert RAM(10398) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10398)))) severity failure;
    assert RAM(10399) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10399)))) severity failure;
    assert RAM(10400) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10400)))) severity failure;
    assert RAM(10401) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10401)))) severity failure;
    assert RAM(10402) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10402)))) severity failure;
    assert RAM(10403) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10403)))) severity failure;
    assert RAM(10404) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10404)))) severity failure;
    assert RAM(10405) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10405)))) severity failure;
    assert RAM(10406) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10406)))) severity failure;
    assert RAM(10407) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10407)))) severity failure;
    assert RAM(10408) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10408)))) severity failure;
    assert RAM(10409) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10409)))) severity failure;
    assert RAM(10410) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10410)))) severity failure;
    assert RAM(10411) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10411)))) severity failure;
    assert RAM(10412) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10412)))) severity failure;
    assert RAM(10413) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10413)))) severity failure;
    assert RAM(10414) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10414)))) severity failure;
    assert RAM(10415) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10415)))) severity failure;
    assert RAM(10416) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10416)))) severity failure;
    assert RAM(10417) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10417)))) severity failure;
    assert RAM(10418) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10418)))) severity failure;
    assert RAM(10419) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10419)))) severity failure;
    assert RAM(10420) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10420)))) severity failure;
    assert RAM(10421) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10421)))) severity failure;
    assert RAM(10422) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10422)))) severity failure;
    assert RAM(10423) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10423)))) severity failure;
    assert RAM(10424) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10424)))) severity failure;
    assert RAM(10425) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10425)))) severity failure;
    assert RAM(10426) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10426)))) severity failure;
    assert RAM(10427) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10427)))) severity failure;
    assert RAM(10428) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10428)))) severity failure;
    assert RAM(10429) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10429)))) severity failure;
    assert RAM(10430) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10430)))) severity failure;
    assert RAM(10431) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10431)))) severity failure;
    assert RAM(10432) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10432)))) severity failure;
    assert RAM(10433) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10433)))) severity failure;
    assert RAM(10434) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10434)))) severity failure;
    assert RAM(10435) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10435)))) severity failure;
    assert RAM(10436) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10436)))) severity failure;
    assert RAM(10437) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10437)))) severity failure;
    assert RAM(10438) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10438)))) severity failure;
    assert RAM(10439) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10439)))) severity failure;
    assert RAM(10440) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10440)))) severity failure;
    assert RAM(10441) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10441)))) severity failure;
    assert RAM(10442) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10442)))) severity failure;
    assert RAM(10443) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10443)))) severity failure;
    assert RAM(10444) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10444)))) severity failure;
    assert RAM(10445) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10445)))) severity failure;
    assert RAM(10446) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10446)))) severity failure;
    assert RAM(10447) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10447)))) severity failure;
    assert RAM(10448) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10448)))) severity failure;
    assert RAM(10449) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10449)))) severity failure;
    assert RAM(10450) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10450)))) severity failure;
    assert RAM(10451) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10451)))) severity failure;
    assert RAM(10452) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10452)))) severity failure;
    assert RAM(10453) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10453)))) severity failure;
    assert RAM(10454) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10454)))) severity failure;
    assert RAM(10455) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10455)))) severity failure;
    assert RAM(10456) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10456)))) severity failure;
    assert RAM(10457) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10457)))) severity failure;
    assert RAM(10458) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10458)))) severity failure;
    assert RAM(10459) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10459)))) severity failure;
    assert RAM(10460) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10460)))) severity failure;
    assert RAM(10461) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10461)))) severity failure;
    assert RAM(10462) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10462)))) severity failure;
    assert RAM(10463) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10463)))) severity failure;
    assert RAM(10464) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10464)))) severity failure;
    assert RAM(10465) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10465)))) severity failure;
    assert RAM(10466) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10466)))) severity failure;
    assert RAM(10467) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10467)))) severity failure;
    assert RAM(10468) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10468)))) severity failure;
    assert RAM(10469) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10469)))) severity failure;
    assert RAM(10470) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10470)))) severity failure;
    assert RAM(10471) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10471)))) severity failure;
    assert RAM(10472) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10472)))) severity failure;
    assert RAM(10473) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10473)))) severity failure;
    assert RAM(10474) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10474)))) severity failure;
    assert RAM(10475) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10475)))) severity failure;
    assert RAM(10476) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10476)))) severity failure;
    assert RAM(10477) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10477)))) severity failure;
    assert RAM(10478) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10478)))) severity failure;
    assert RAM(10479) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10479)))) severity failure;
    assert RAM(10480) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10480)))) severity failure;
    assert RAM(10481) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10481)))) severity failure;
    assert RAM(10482) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10482)))) severity failure;
    assert RAM(10483) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10483)))) severity failure;
    assert RAM(10484) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10484)))) severity failure;
    assert RAM(10485) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10485)))) severity failure;
    assert RAM(10486) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10486)))) severity failure;
    assert RAM(10487) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10487)))) severity failure;
    assert RAM(10488) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10488)))) severity failure;
    assert RAM(10489) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10489)))) severity failure;
    assert RAM(10490) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10490)))) severity failure;
    assert RAM(10491) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10491)))) severity failure;
    assert RAM(10492) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10492)))) severity failure;
    assert RAM(10493) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10493)))) severity failure;
    assert RAM(10494) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10494)))) severity failure;
    assert RAM(10495) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10495)))) severity failure;
    assert RAM(10496) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10496)))) severity failure;
    assert RAM(10497) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10497)))) severity failure;
    assert RAM(10498) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10498)))) severity failure;
    assert RAM(10499) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10499)))) severity failure;
    assert RAM(10500) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10500)))) severity failure;
    assert RAM(10501) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10501)))) severity failure;
    assert RAM(10502) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10502)))) severity failure;
    assert RAM(10503) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10503)))) severity failure;
    assert RAM(10504) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10504)))) severity failure;
    assert RAM(10505) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10505)))) severity failure;
    assert RAM(10506) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10506)))) severity failure;
    assert RAM(10507) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10507)))) severity failure;
    assert RAM(10508) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10508)))) severity failure;
    assert RAM(10509) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10509)))) severity failure;
    assert RAM(10510) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10510)))) severity failure;
    assert RAM(10511) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10511)))) severity failure;
    assert RAM(10512) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10512)))) severity failure;
    assert RAM(10513) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10513)))) severity failure;
    assert RAM(10514) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10514)))) severity failure;
    assert RAM(10515) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10515)))) severity failure;
    assert RAM(10516) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10516)))) severity failure;
    assert RAM(10517) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10517)))) severity failure;
    assert RAM(10518) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10518)))) severity failure;
    assert RAM(10519) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10519)))) severity failure;
    assert RAM(10520) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10520)))) severity failure;
    assert RAM(10521) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10521)))) severity failure;
    assert RAM(10522) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10522)))) severity failure;
    assert RAM(10523) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10523)))) severity failure;
    assert RAM(10524) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10524)))) severity failure;
    assert RAM(10525) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10525)))) severity failure;
    assert RAM(10526) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10526)))) severity failure;
    assert RAM(10527) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10527)))) severity failure;
    assert RAM(10528) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10528)))) severity failure;
    assert RAM(10529) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10529)))) severity failure;
    assert RAM(10530) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10530)))) severity failure;
    assert RAM(10531) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10531)))) severity failure;
    assert RAM(10532) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10532)))) severity failure;
    assert RAM(10533) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10533)))) severity failure;
    assert RAM(10534) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10534)))) severity failure;
    assert RAM(10535) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10535)))) severity failure;
    assert RAM(10536) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10536)))) severity failure;
    assert RAM(10537) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10537)))) severity failure;
    assert RAM(10538) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10538)))) severity failure;
    assert RAM(10539) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10539)))) severity failure;
    assert RAM(10540) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10540)))) severity failure;
    assert RAM(10541) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10541)))) severity failure;
    assert RAM(10542) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10542)))) severity failure;
    assert RAM(10543) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10543)))) severity failure;
    assert RAM(10544) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10544)))) severity failure;
    assert RAM(10545) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10545)))) severity failure;
    assert RAM(10546) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10546)))) severity failure;
    assert RAM(10547) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10547)))) severity failure;
    assert RAM(10548) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10548)))) severity failure;
    assert RAM(10549) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10549)))) severity failure;
    assert RAM(10550) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10550)))) severity failure;
    assert RAM(10551) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10551)))) severity failure;
    assert RAM(10552) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10552)))) severity failure;
    assert RAM(10553) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10553)))) severity failure;
    assert RAM(10554) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10554)))) severity failure;
    assert RAM(10555) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10555)))) severity failure;
    assert RAM(10556) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10556)))) severity failure;
    assert RAM(10557) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10557)))) severity failure;
    assert RAM(10558) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10558)))) severity failure;
    assert RAM(10559) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10559)))) severity failure;
    assert RAM(10560) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10560)))) severity failure;
    assert RAM(10561) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10561)))) severity failure;
    assert RAM(10562) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10562)))) severity failure;
    assert RAM(10563) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10563)))) severity failure;
    assert RAM(10564) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10564)))) severity failure;
    assert RAM(10565) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10565)))) severity failure;
    assert RAM(10566) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10566)))) severity failure;
    assert RAM(10567) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10567)))) severity failure;
    assert RAM(10568) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10568)))) severity failure;
    assert RAM(10569) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10569)))) severity failure;
    assert RAM(10570) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10570)))) severity failure;
    assert RAM(10571) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10571)))) severity failure;
    assert RAM(10572) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10572)))) severity failure;
    assert RAM(10573) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10573)))) severity failure;
    assert RAM(10574) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10574)))) severity failure;
    assert RAM(10575) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10575)))) severity failure;
    assert RAM(10576) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10576)))) severity failure;
    assert RAM(10577) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10577)))) severity failure;
    assert RAM(10578) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10578)))) severity failure;
    assert RAM(10579) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10579)))) severity failure;
    assert RAM(10580) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10580)))) severity failure;
    assert RAM(10581) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10581)))) severity failure;
    assert RAM(10582) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10582)))) severity failure;
    assert RAM(10583) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10583)))) severity failure;
    assert RAM(10584) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10584)))) severity failure;
    assert RAM(10585) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10585)))) severity failure;
    assert RAM(10586) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10586)))) severity failure;
    assert RAM(10587) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10587)))) severity failure;
    assert RAM(10588) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10588)))) severity failure;
    assert RAM(10589) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10589)))) severity failure;
    assert RAM(10590) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10590)))) severity failure;
    assert RAM(10591) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10591)))) severity failure;
    assert RAM(10592) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10592)))) severity failure;
    assert RAM(10593) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10593)))) severity failure;
    assert RAM(10594) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10594)))) severity failure;
    assert RAM(10595) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10595)))) severity failure;
    assert RAM(10596) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10596)))) severity failure;
    assert RAM(10597) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10597)))) severity failure;
    assert RAM(10598) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10598)))) severity failure;
    assert RAM(10599) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10599)))) severity failure;
    assert RAM(10600) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10600)))) severity failure;
    assert RAM(10601) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10601)))) severity failure;
    assert RAM(10602) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10602)))) severity failure;
    assert RAM(10603) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10603)))) severity failure;
    assert RAM(10604) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10604)))) severity failure;
    assert RAM(10605) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10605)))) severity failure;
    assert RAM(10606) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10606)))) severity failure;
    assert RAM(10607) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10607)))) severity failure;
    assert RAM(10608) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10608)))) severity failure;
    assert RAM(10609) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10609)))) severity failure;
    assert RAM(10610) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10610)))) severity failure;
    assert RAM(10611) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10611)))) severity failure;
    assert RAM(10612) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10612)))) severity failure;
    assert RAM(10613) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10613)))) severity failure;
    assert RAM(10614) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10614)))) severity failure;
    assert RAM(10615) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10615)))) severity failure;
    assert RAM(10616) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10616)))) severity failure;
    assert RAM(10617) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10617)))) severity failure;
    assert RAM(10618) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10618)))) severity failure;
    assert RAM(10619) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10619)))) severity failure;
    assert RAM(10620) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10620)))) severity failure;
    assert RAM(10621) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10621)))) severity failure;
    assert RAM(10622) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10622)))) severity failure;
    assert RAM(10623) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10623)))) severity failure;
    assert RAM(10624) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10624)))) severity failure;
    assert RAM(10625) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10625)))) severity failure;
    assert RAM(10626) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10626)))) severity failure;
    assert RAM(10627) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10627)))) severity failure;
    assert RAM(10628) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10628)))) severity failure;
    assert RAM(10629) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10629)))) severity failure;
    assert RAM(10630) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10630)))) severity failure;
    assert RAM(10631) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10631)))) severity failure;
    assert RAM(10632) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10632)))) severity failure;
    assert RAM(10633) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10633)))) severity failure;
    assert RAM(10634) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10634)))) severity failure;
    assert RAM(10635) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10635)))) severity failure;
    assert RAM(10636) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10636)))) severity failure;
    assert RAM(10637) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10637)))) severity failure;
    assert RAM(10638) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10638)))) severity failure;
    assert RAM(10639) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10639)))) severity failure;
    assert RAM(10640) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10640)))) severity failure;
    assert RAM(10641) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10641)))) severity failure;
    assert RAM(10642) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10642)))) severity failure;
    assert RAM(10643) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10643)))) severity failure;
    assert RAM(10644) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10644)))) severity failure;
    assert RAM(10645) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10645)))) severity failure;
    assert RAM(10646) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10646)))) severity failure;
    assert RAM(10647) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10647)))) severity failure;
    assert RAM(10648) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10648)))) severity failure;
    assert RAM(10649) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10649)))) severity failure;
    assert RAM(10650) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10650)))) severity failure;
    assert RAM(10651) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10651)))) severity failure;
    assert RAM(10652) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10652)))) severity failure;
    assert RAM(10653) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10653)))) severity failure;
    assert RAM(10654) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10654)))) severity failure;
    assert RAM(10655) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10655)))) severity failure;
    assert RAM(10656) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10656)))) severity failure;
    assert RAM(10657) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10657)))) severity failure;
    assert RAM(10658) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10658)))) severity failure;
    assert RAM(10659) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10659)))) severity failure;
    assert RAM(10660) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10660)))) severity failure;
    assert RAM(10661) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10661)))) severity failure;
    assert RAM(10662) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10662)))) severity failure;
    assert RAM(10663) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10663)))) severity failure;
    assert RAM(10664) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10664)))) severity failure;
    assert RAM(10665) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10665)))) severity failure;
    assert RAM(10666) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10666)))) severity failure;
    assert RAM(10667) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10667)))) severity failure;
    assert RAM(10668) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10668)))) severity failure;
    assert RAM(10669) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10669)))) severity failure;
    assert RAM(10670) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10670)))) severity failure;
    assert RAM(10671) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10671)))) severity failure;
    assert RAM(10672) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10672)))) severity failure;
    assert RAM(10673) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10673)))) severity failure;
    assert RAM(10674) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10674)))) severity failure;
    assert RAM(10675) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10675)))) severity failure;
    assert RAM(10676) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10676)))) severity failure;
    assert RAM(10677) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10677)))) severity failure;
    assert RAM(10678) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10678)))) severity failure;
    assert RAM(10679) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10679)))) severity failure;
    assert RAM(10680) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10680)))) severity failure;
    assert RAM(10681) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10681)))) severity failure;
    assert RAM(10682) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10682)))) severity failure;
    assert RAM(10683) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10683)))) severity failure;
    assert RAM(10684) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10684)))) severity failure;
    assert RAM(10685) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10685)))) severity failure;
    assert RAM(10686) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10686)))) severity failure;
    assert RAM(10687) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10687)))) severity failure;
    assert RAM(10688) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10688)))) severity failure;
    assert RAM(10689) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10689)))) severity failure;
    assert RAM(10690) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10690)))) severity failure;
    assert RAM(10691) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10691)))) severity failure;
    assert RAM(10692) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10692)))) severity failure;
    assert RAM(10693) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10693)))) severity failure;
    assert RAM(10694) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10694)))) severity failure;
    assert RAM(10695) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10695)))) severity failure;
    assert RAM(10696) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10696)))) severity failure;
    assert RAM(10697) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10697)))) severity failure;
    assert RAM(10698) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10698)))) severity failure;
    assert RAM(10699) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10699)))) severity failure;
    assert RAM(10700) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10700)))) severity failure;
    assert RAM(10701) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10701)))) severity failure;
    assert RAM(10702) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10702)))) severity failure;
    assert RAM(10703) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10703)))) severity failure;
    assert RAM(10704) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10704)))) severity failure;
    assert RAM(10705) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10705)))) severity failure;
    assert RAM(10706) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10706)))) severity failure;
    assert RAM(10707) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10707)))) severity failure;
    assert RAM(10708) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10708)))) severity failure;
    assert RAM(10709) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10709)))) severity failure;
    assert RAM(10710) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10710)))) severity failure;
    assert RAM(10711) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10711)))) severity failure;
    assert RAM(10712) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10712)))) severity failure;
    assert RAM(10713) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10713)))) severity failure;
    assert RAM(10714) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10714)))) severity failure;
    assert RAM(10715) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10715)))) severity failure;
    assert RAM(10716) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10716)))) severity failure;
    assert RAM(10717) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10717)))) severity failure;
    assert RAM(10718) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10718)))) severity failure;
    assert RAM(10719) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10719)))) severity failure;
    assert RAM(10720) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10720)))) severity failure;
    assert RAM(10721) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10721)))) severity failure;
    assert RAM(10722) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10722)))) severity failure;
    assert RAM(10723) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10723)))) severity failure;
    assert RAM(10724) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10724)))) severity failure;
    assert RAM(10725) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10725)))) severity failure;
    assert RAM(10726) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10726)))) severity failure;
    assert RAM(10727) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10727)))) severity failure;
    assert RAM(10728) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10728)))) severity failure;
    assert RAM(10729) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10729)))) severity failure;
    assert RAM(10730) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10730)))) severity failure;
    assert RAM(10731) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10731)))) severity failure;
    assert RAM(10732) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10732)))) severity failure;
    assert RAM(10733) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10733)))) severity failure;
    assert RAM(10734) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10734)))) severity failure;
    assert RAM(10735) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10735)))) severity failure;
    assert RAM(10736) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10736)))) severity failure;
    assert RAM(10737) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10737)))) severity failure;
    assert RAM(10738) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10738)))) severity failure;
    assert RAM(10739) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10739)))) severity failure;
    assert RAM(10740) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10740)))) severity failure;
    assert RAM(10741) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10741)))) severity failure;
    assert RAM(10742) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10742)))) severity failure;
    assert RAM(10743) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10743)))) severity failure;
    assert RAM(10744) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10744)))) severity failure;
    assert RAM(10745) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10745)))) severity failure;
    assert RAM(10746) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10746)))) severity failure;
    assert RAM(10747) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10747)))) severity failure;
    assert RAM(10748) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10748)))) severity failure;
    assert RAM(10749) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10749)))) severity failure;
    assert RAM(10750) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10750)))) severity failure;
    assert RAM(10751) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10751)))) severity failure;
    assert RAM(10752) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10752)))) severity failure;
    assert RAM(10753) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10753)))) severity failure;
    assert RAM(10754) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10754)))) severity failure;
    assert RAM(10755) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10755)))) severity failure;
    assert RAM(10756) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10756)))) severity failure;
    assert RAM(10757) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10757)))) severity failure;
    assert RAM(10758) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10758)))) severity failure;
    assert RAM(10759) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10759)))) severity failure;
    assert RAM(10760) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10760)))) severity failure;
    assert RAM(10761) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10761)))) severity failure;
    assert RAM(10762) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10762)))) severity failure;
    assert RAM(10763) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10763)))) severity failure;
    assert RAM(10764) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10764)))) severity failure;
    assert RAM(10765) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10765)))) severity failure;
    assert RAM(10766) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10766)))) severity failure;
    assert RAM(10767) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10767)))) severity failure;
    assert RAM(10768) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10768)))) severity failure;
    assert RAM(10769) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10769)))) severity failure;
    assert RAM(10770) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10770)))) severity failure;
    assert RAM(10771) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10771)))) severity failure;
    assert RAM(10772) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10772)))) severity failure;
    assert RAM(10773) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10773)))) severity failure;
    assert RAM(10774) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10774)))) severity failure;
    assert RAM(10775) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10775)))) severity failure;
    assert RAM(10776) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10776)))) severity failure;
    assert RAM(10777) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10777)))) severity failure;
    assert RAM(10778) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10778)))) severity failure;
    assert RAM(10779) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10779)))) severity failure;
    assert RAM(10780) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10780)))) severity failure;
    assert RAM(10781) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10781)))) severity failure;
    assert RAM(10782) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10782)))) severity failure;
    assert RAM(10783) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10783)))) severity failure;
    assert RAM(10784) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10784)))) severity failure;
    assert RAM(10785) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10785)))) severity failure;
    assert RAM(10786) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10786)))) severity failure;
    assert RAM(10787) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10787)))) severity failure;
    assert RAM(10788) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10788)))) severity failure;
    assert RAM(10789) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10789)))) severity failure;
    assert RAM(10790) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10790)))) severity failure;
    assert RAM(10791) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10791)))) severity failure;
    assert RAM(10792) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10792)))) severity failure;
    assert RAM(10793) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10793)))) severity failure;
    assert RAM(10794) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10794)))) severity failure;
    assert RAM(10795) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10795)))) severity failure;
    assert RAM(10796) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10796)))) severity failure;
    assert RAM(10797) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10797)))) severity failure;
    assert RAM(10798) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10798)))) severity failure;
    assert RAM(10799) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10799)))) severity failure;
    assert RAM(10800) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10800)))) severity failure;
    assert RAM(10801) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10801)))) severity failure;
    assert RAM(10802) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10802)))) severity failure;
    assert RAM(10803) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10803)))) severity failure;
    assert RAM(10804) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10804)))) severity failure;
    assert RAM(10805) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10805)))) severity failure;
    assert RAM(10806) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10806)))) severity failure;
    assert RAM(10807) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10807)))) severity failure;
    assert RAM(10808) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10808)))) severity failure;
    assert RAM(10809) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10809)))) severity failure;
    assert RAM(10810) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10810)))) severity failure;
    assert RAM(10811) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10811)))) severity failure;
    assert RAM(10812) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10812)))) severity failure;
    assert RAM(10813) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10813)))) severity failure;
    assert RAM(10814) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10814)))) severity failure;
    assert RAM(10815) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10815)))) severity failure;
    assert RAM(10816) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10816)))) severity failure;
    assert RAM(10817) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10817)))) severity failure;
    assert RAM(10818) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10818)))) severity failure;
    assert RAM(10819) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10819)))) severity failure;
    assert RAM(10820) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10820)))) severity failure;
    assert RAM(10821) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10821)))) severity failure;
    assert RAM(10822) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10822)))) severity failure;
    assert RAM(10823) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10823)))) severity failure;
    assert RAM(10824) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10824)))) severity failure;
    assert RAM(10825) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10825)))) severity failure;
    assert RAM(10826) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10826)))) severity failure;
    assert RAM(10827) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10827)))) severity failure;
    assert RAM(10828) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10828)))) severity failure;
    assert RAM(10829) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10829)))) severity failure;
    assert RAM(10830) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10830)))) severity failure;
    assert RAM(10831) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10831)))) severity failure;
    assert RAM(10832) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10832)))) severity failure;
    assert RAM(10833) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10833)))) severity failure;
    assert RAM(10834) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10834)))) severity failure;
    assert RAM(10835) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10835)))) severity failure;
    assert RAM(10836) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10836)))) severity failure;
    assert RAM(10837) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10837)))) severity failure;
    assert RAM(10838) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10838)))) severity failure;
    assert RAM(10839) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10839)))) severity failure;
    assert RAM(10840) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10840)))) severity failure;
    assert RAM(10841) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10841)))) severity failure;
    assert RAM(10842) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10842)))) severity failure;
    assert RAM(10843) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10843)))) severity failure;
    assert RAM(10844) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10844)))) severity failure;
    assert RAM(10845) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10845)))) severity failure;
    assert RAM(10846) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10846)))) severity failure;
    assert RAM(10847) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10847)))) severity failure;
    assert RAM(10848) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10848)))) severity failure;
    assert RAM(10849) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10849)))) severity failure;
    assert RAM(10850) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10850)))) severity failure;
    assert RAM(10851) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10851)))) severity failure;
    assert RAM(10852) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10852)))) severity failure;
    assert RAM(10853) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10853)))) severity failure;
    assert RAM(10854) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10854)))) severity failure;
    assert RAM(10855) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10855)))) severity failure;
    assert RAM(10856) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10856)))) severity failure;
    assert RAM(10857) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10857)))) severity failure;
    assert RAM(10858) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10858)))) severity failure;
    assert RAM(10859) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10859)))) severity failure;
    assert RAM(10860) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10860)))) severity failure;
    assert RAM(10861) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10861)))) severity failure;
    assert RAM(10862) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10862)))) severity failure;
    assert RAM(10863) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10863)))) severity failure;
    assert RAM(10864) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10864)))) severity failure;
    assert RAM(10865) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10865)))) severity failure;
    assert RAM(10866) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10866)))) severity failure;
    assert RAM(10867) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10867)))) severity failure;
    assert RAM(10868) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10868)))) severity failure;
    assert RAM(10869) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10869)))) severity failure;
    assert RAM(10870) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10870)))) severity failure;
    assert RAM(10871) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10871)))) severity failure;
    assert RAM(10872) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10872)))) severity failure;
    assert RAM(10873) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10873)))) severity failure;
    assert RAM(10874) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10874)))) severity failure;
    assert RAM(10875) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10875)))) severity failure;
    assert RAM(10876) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10876)))) severity failure;
    assert RAM(10877) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10877)))) severity failure;
    assert RAM(10878) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10878)))) severity failure;
    assert RAM(10879) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10879)))) severity failure;
    assert RAM(10880) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10880)))) severity failure;
    assert RAM(10881) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10881)))) severity failure;
    assert RAM(10882) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10882)))) severity failure;
    assert RAM(10883) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10883)))) severity failure;
    assert RAM(10884) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10884)))) severity failure;
    assert RAM(10885) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10885)))) severity failure;
    assert RAM(10886) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10886)))) severity failure;
    assert RAM(10887) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10887)))) severity failure;
    assert RAM(10888) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10888)))) severity failure;
    assert RAM(10889) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10889)))) severity failure;
    assert RAM(10890) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10890)))) severity failure;
    assert RAM(10891) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10891)))) severity failure;
    assert RAM(10892) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10892)))) severity failure;
    assert RAM(10893) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10893)))) severity failure;
    assert RAM(10894) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10894)))) severity failure;
    assert RAM(10895) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10895)))) severity failure;
    assert RAM(10896) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10896)))) severity failure;
    assert RAM(10897) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10897)))) severity failure;
    assert RAM(10898) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10898)))) severity failure;
    assert RAM(10899) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10899)))) severity failure;
    assert RAM(10900) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10900)))) severity failure;
    assert RAM(10901) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10901)))) severity failure;
    assert RAM(10902) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10902)))) severity failure;
    assert RAM(10903) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10903)))) severity failure;
    assert RAM(10904) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10904)))) severity failure;
    assert RAM(10905) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10905)))) severity failure;
    assert RAM(10906) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10906)))) severity failure;
    assert RAM(10907) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10907)))) severity failure;
    assert RAM(10908) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10908)))) severity failure;
    assert RAM(10909) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10909)))) severity failure;
    assert RAM(10910) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10910)))) severity failure;
    assert RAM(10911) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10911)))) severity failure;
    assert RAM(10912) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10912)))) severity failure;
    assert RAM(10913) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10913)))) severity failure;
    assert RAM(10914) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10914)))) severity failure;
    assert RAM(10915) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10915)))) severity failure;
    assert RAM(10916) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10916)))) severity failure;
    assert RAM(10917) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10917)))) severity failure;
    assert RAM(10918) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10918)))) severity failure;
    assert RAM(10919) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10919)))) severity failure;
    assert RAM(10920) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10920)))) severity failure;
    assert RAM(10921) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10921)))) severity failure;
    assert RAM(10922) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10922)))) severity failure;
    assert RAM(10923) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10923)))) severity failure;
    assert RAM(10924) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10924)))) severity failure;
    assert RAM(10925) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10925)))) severity failure;
    assert RAM(10926) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10926)))) severity failure;
    assert RAM(10927) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10927)))) severity failure;
    assert RAM(10928) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10928)))) severity failure;
    assert RAM(10929) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10929)))) severity failure;
    assert RAM(10930) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10930)))) severity failure;
    assert RAM(10931) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10931)))) severity failure;
    assert RAM(10932) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10932)))) severity failure;
    assert RAM(10933) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10933)))) severity failure;
    assert RAM(10934) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10934)))) severity failure;
    assert RAM(10935) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10935)))) severity failure;
    assert RAM(10936) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10936)))) severity failure;
    assert RAM(10937) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10937)))) severity failure;
    assert RAM(10938) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10938)))) severity failure;
    assert RAM(10939) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10939)))) severity failure;
    assert RAM(10940) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10940)))) severity failure;
    assert RAM(10941) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10941)))) severity failure;
    assert RAM(10942) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10942)))) severity failure;
    assert RAM(10943) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10943)))) severity failure;
    assert RAM(10944) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10944)))) severity failure;
    assert RAM(10945) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10945)))) severity failure;
    assert RAM(10946) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10946)))) severity failure;
    assert RAM(10947) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10947)))) severity failure;
    assert RAM(10948) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10948)))) severity failure;
    assert RAM(10949) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10949)))) severity failure;
    assert RAM(10950) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10950)))) severity failure;
    assert RAM(10951) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10951)))) severity failure;
    assert RAM(10952) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10952)))) severity failure;
    assert RAM(10953) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10953)))) severity failure;
    assert RAM(10954) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10954)))) severity failure;
    assert RAM(10955) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10955)))) severity failure;
    assert RAM(10956) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10956)))) severity failure;
    assert RAM(10957) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10957)))) severity failure;
    assert RAM(10958) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10958)))) severity failure;
    assert RAM(10959) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10959)))) severity failure;
    assert RAM(10960) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10960)))) severity failure;
    assert RAM(10961) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10961)))) severity failure;
    assert RAM(10962) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10962)))) severity failure;
    assert RAM(10963) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10963)))) severity failure;
    assert RAM(10964) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10964)))) severity failure;
    assert RAM(10965) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10965)))) severity failure;
    assert RAM(10966) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10966)))) severity failure;
    assert RAM(10967) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10967)))) severity failure;
    assert RAM(10968) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10968)))) severity failure;
    assert RAM(10969) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10969)))) severity failure;
    assert RAM(10970) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10970)))) severity failure;
    assert RAM(10971) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10971)))) severity failure;
    assert RAM(10972) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10972)))) severity failure;
    assert RAM(10973) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10973)))) severity failure;
    assert RAM(10974) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10974)))) severity failure;
    assert RAM(10975) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10975)))) severity failure;
    assert RAM(10976) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10976)))) severity failure;
    assert RAM(10977) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10977)))) severity failure;
    assert RAM(10978) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10978)))) severity failure;
    assert RAM(10979) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10979)))) severity failure;
    assert RAM(10980) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10980)))) severity failure;
    assert RAM(10981) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10981)))) severity failure;
    assert RAM(10982) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10982)))) severity failure;
    assert RAM(10983) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10983)))) severity failure;
    assert RAM(10984) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10984)))) severity failure;
    assert RAM(10985) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10985)))) severity failure;
    assert RAM(10986) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10986)))) severity failure;
    assert RAM(10987) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10987)))) severity failure;
    assert RAM(10988) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10988)))) severity failure;
    assert RAM(10989) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10989)))) severity failure;
    assert RAM(10990) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10990)))) severity failure;
    assert RAM(10991) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10991)))) severity failure;
    assert RAM(10992) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10992)))) severity failure;
    assert RAM(10993) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10993)))) severity failure;
    assert RAM(10994) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10994)))) severity failure;
    assert RAM(10995) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10995)))) severity failure;
    assert RAM(10996) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10996)))) severity failure;
    assert RAM(10997) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(10997)))) severity failure;
    assert RAM(10998) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10998)))) severity failure;
    assert RAM(10999) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(10999)))) severity failure;
    assert RAM(11000) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11000)))) severity failure;
    assert RAM(11001) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11001)))) severity failure;
    assert RAM(11002) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11002)))) severity failure;
    assert RAM(11003) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11003)))) severity failure;
    assert RAM(11004) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11004)))) severity failure;
    assert RAM(11005) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11005)))) severity failure;
    assert RAM(11006) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11006)))) severity failure;
    assert RAM(11007) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11007)))) severity failure;
    assert RAM(11008) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11008)))) severity failure;
    assert RAM(11009) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11009)))) severity failure;
    assert RAM(11010) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11010)))) severity failure;
    assert RAM(11011) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11011)))) severity failure;
    assert RAM(11012) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11012)))) severity failure;
    assert RAM(11013) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11013)))) severity failure;
    assert RAM(11014) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11014)))) severity failure;
    assert RAM(11015) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11015)))) severity failure;
    assert RAM(11016) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11016)))) severity failure;
    assert RAM(11017) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11017)))) severity failure;
    assert RAM(11018) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11018)))) severity failure;
    assert RAM(11019) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11019)))) severity failure;
    assert RAM(11020) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11020)))) severity failure;
    assert RAM(11021) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11021)))) severity failure;
    assert RAM(11022) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11022)))) severity failure;
    assert RAM(11023) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11023)))) severity failure;
    assert RAM(11024) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11024)))) severity failure;
    assert RAM(11025) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11025)))) severity failure;
    assert RAM(11026) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11026)))) severity failure;
    assert RAM(11027) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11027)))) severity failure;
    assert RAM(11028) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11028)))) severity failure;
    assert RAM(11029) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11029)))) severity failure;
    assert RAM(11030) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11030)))) severity failure;
    assert RAM(11031) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11031)))) severity failure;
    assert RAM(11032) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11032)))) severity failure;
    assert RAM(11033) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11033)))) severity failure;
    assert RAM(11034) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11034)))) severity failure;
    assert RAM(11035) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11035)))) severity failure;
    assert RAM(11036) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11036)))) severity failure;
    assert RAM(11037) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11037)))) severity failure;
    assert RAM(11038) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11038)))) severity failure;
    assert RAM(11039) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11039)))) severity failure;
    assert RAM(11040) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11040)))) severity failure;
    assert RAM(11041) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11041)))) severity failure;
    assert RAM(11042) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11042)))) severity failure;
    assert RAM(11043) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11043)))) severity failure;
    assert RAM(11044) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11044)))) severity failure;
    assert RAM(11045) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11045)))) severity failure;
    assert RAM(11046) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11046)))) severity failure;
    assert RAM(11047) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11047)))) severity failure;
    assert RAM(11048) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11048)))) severity failure;
    assert RAM(11049) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11049)))) severity failure;
    assert RAM(11050) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11050)))) severity failure;
    assert RAM(11051) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11051)))) severity failure;
    assert RAM(11052) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11052)))) severity failure;
    assert RAM(11053) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11053)))) severity failure;
    assert RAM(11054) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11054)))) severity failure;
    assert RAM(11055) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11055)))) severity failure;
    assert RAM(11056) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11056)))) severity failure;
    assert RAM(11057) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11057)))) severity failure;
    assert RAM(11058) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11058)))) severity failure;
    assert RAM(11059) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11059)))) severity failure;
    assert RAM(11060) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11060)))) severity failure;
    assert RAM(11061) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11061)))) severity failure;
    assert RAM(11062) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11062)))) severity failure;
    assert RAM(11063) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11063)))) severity failure;
    assert RAM(11064) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11064)))) severity failure;
    assert RAM(11065) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11065)))) severity failure;
    assert RAM(11066) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11066)))) severity failure;
    assert RAM(11067) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11067)))) severity failure;
    assert RAM(11068) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11068)))) severity failure;
    assert RAM(11069) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11069)))) severity failure;
    assert RAM(11070) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11070)))) severity failure;
    assert RAM(11071) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11071)))) severity failure;
    assert RAM(11072) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11072)))) severity failure;
    assert RAM(11073) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11073)))) severity failure;
    assert RAM(11074) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11074)))) severity failure;
    assert RAM(11075) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11075)))) severity failure;
    assert RAM(11076) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11076)))) severity failure;
    assert RAM(11077) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11077)))) severity failure;
    assert RAM(11078) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11078)))) severity failure;
    assert RAM(11079) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11079)))) severity failure;
    assert RAM(11080) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11080)))) severity failure;
    assert RAM(11081) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11081)))) severity failure;
    assert RAM(11082) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11082)))) severity failure;
    assert RAM(11083) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11083)))) severity failure;
    assert RAM(11084) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11084)))) severity failure;
    assert RAM(11085) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11085)))) severity failure;
    assert RAM(11086) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11086)))) severity failure;
    assert RAM(11087) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11087)))) severity failure;
    assert RAM(11088) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11088)))) severity failure;
    assert RAM(11089) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11089)))) severity failure;
    assert RAM(11090) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11090)))) severity failure;
    assert RAM(11091) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11091)))) severity failure;
    assert RAM(11092) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11092)))) severity failure;
    assert RAM(11093) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11093)))) severity failure;
    assert RAM(11094) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11094)))) severity failure;
    assert RAM(11095) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11095)))) severity failure;
    assert RAM(11096) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11096)))) severity failure;
    assert RAM(11097) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11097)))) severity failure;
    assert RAM(11098) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11098)))) severity failure;
    assert RAM(11099) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11099)))) severity failure;
    assert RAM(11100) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11100)))) severity failure;
    assert RAM(11101) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11101)))) severity failure;
    assert RAM(11102) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11102)))) severity failure;
    assert RAM(11103) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11103)))) severity failure;
    assert RAM(11104) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11104)))) severity failure;
    assert RAM(11105) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11105)))) severity failure;
    assert RAM(11106) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11106)))) severity failure;
    assert RAM(11107) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11107)))) severity failure;
    assert RAM(11108) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11108)))) severity failure;
    assert RAM(11109) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11109)))) severity failure;
    assert RAM(11110) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11110)))) severity failure;
    assert RAM(11111) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11111)))) severity failure;
    assert RAM(11112) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11112)))) severity failure;
    assert RAM(11113) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11113)))) severity failure;
    assert RAM(11114) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11114)))) severity failure;
    assert RAM(11115) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11115)))) severity failure;
    assert RAM(11116) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11116)))) severity failure;
    assert RAM(11117) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11117)))) severity failure;
    assert RAM(11118) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11118)))) severity failure;
    assert RAM(11119) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11119)))) severity failure;
    assert RAM(11120) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11120)))) severity failure;
    assert RAM(11121) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11121)))) severity failure;
    assert RAM(11122) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11122)))) severity failure;
    assert RAM(11123) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11123)))) severity failure;
    assert RAM(11124) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11124)))) severity failure;
    assert RAM(11125) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11125)))) severity failure;
    assert RAM(11126) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11126)))) severity failure;
    assert RAM(11127) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11127)))) severity failure;
    assert RAM(11128) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11128)))) severity failure;
    assert RAM(11129) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11129)))) severity failure;
    assert RAM(11130) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11130)))) severity failure;
    assert RAM(11131) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11131)))) severity failure;
    assert RAM(11132) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11132)))) severity failure;
    assert RAM(11133) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11133)))) severity failure;
    assert RAM(11134) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11134)))) severity failure;
    assert RAM(11135) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11135)))) severity failure;
    assert RAM(11136) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11136)))) severity failure;
    assert RAM(11137) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11137)))) severity failure;
    assert RAM(11138) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11138)))) severity failure;
    assert RAM(11139) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11139)))) severity failure;
    assert RAM(11140) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11140)))) severity failure;
    assert RAM(11141) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11141)))) severity failure;
    assert RAM(11142) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11142)))) severity failure;
    assert RAM(11143) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11143)))) severity failure;
    assert RAM(11144) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11144)))) severity failure;
    assert RAM(11145) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11145)))) severity failure;
    assert RAM(11146) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11146)))) severity failure;
    assert RAM(11147) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11147)))) severity failure;
    assert RAM(11148) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11148)))) severity failure;
    assert RAM(11149) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11149)))) severity failure;
    assert RAM(11150) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11150)))) severity failure;
    assert RAM(11151) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11151)))) severity failure;
    assert RAM(11152) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11152)))) severity failure;
    assert RAM(11153) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11153)))) severity failure;
    assert RAM(11154) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11154)))) severity failure;
    assert RAM(11155) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11155)))) severity failure;
    assert RAM(11156) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11156)))) severity failure;
    assert RAM(11157) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11157)))) severity failure;
    assert RAM(11158) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11158)))) severity failure;
    assert RAM(11159) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11159)))) severity failure;
    assert RAM(11160) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11160)))) severity failure;
    assert RAM(11161) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11161)))) severity failure;
    assert RAM(11162) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11162)))) severity failure;
    assert RAM(11163) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11163)))) severity failure;
    assert RAM(11164) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11164)))) severity failure;
    assert RAM(11165) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11165)))) severity failure;
    assert RAM(11166) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11166)))) severity failure;
    assert RAM(11167) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11167)))) severity failure;
    assert RAM(11168) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11168)))) severity failure;
    assert RAM(11169) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11169)))) severity failure;
    assert RAM(11170) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11170)))) severity failure;
    assert RAM(11171) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11171)))) severity failure;
    assert RAM(11172) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11172)))) severity failure;
    assert RAM(11173) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11173)))) severity failure;
    assert RAM(11174) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11174)))) severity failure;
    assert RAM(11175) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11175)))) severity failure;
    assert RAM(11176) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11176)))) severity failure;
    assert RAM(11177) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11177)))) severity failure;
    assert RAM(11178) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11178)))) severity failure;
    assert RAM(11179) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11179)))) severity failure;
    assert RAM(11180) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11180)))) severity failure;
    assert RAM(11181) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11181)))) severity failure;
    assert RAM(11182) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11182)))) severity failure;
    assert RAM(11183) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11183)))) severity failure;
    assert RAM(11184) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11184)))) severity failure;
    assert RAM(11185) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11185)))) severity failure;
    assert RAM(11186) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11186)))) severity failure;
    assert RAM(11187) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11187)))) severity failure;
    assert RAM(11188) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11188)))) severity failure;
    assert RAM(11189) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11189)))) severity failure;
    assert RAM(11190) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11190)))) severity failure;
    assert RAM(11191) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11191)))) severity failure;
    assert RAM(11192) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11192)))) severity failure;
    assert RAM(11193) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11193)))) severity failure;
    assert RAM(11194) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11194)))) severity failure;
    assert RAM(11195) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11195)))) severity failure;
    assert RAM(11196) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11196)))) severity failure;
    assert RAM(11197) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11197)))) severity failure;
    assert RAM(11198) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11198)))) severity failure;
    assert RAM(11199) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11199)))) severity failure;
    assert RAM(11200) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11200)))) severity failure;
    assert RAM(11201) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11201)))) severity failure;
    assert RAM(11202) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11202)))) severity failure;
    assert RAM(11203) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11203)))) severity failure;
    assert RAM(11204) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11204)))) severity failure;
    assert RAM(11205) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11205)))) severity failure;
    assert RAM(11206) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11206)))) severity failure;
    assert RAM(11207) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11207)))) severity failure;
    assert RAM(11208) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11208)))) severity failure;
    assert RAM(11209) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11209)))) severity failure;
    assert RAM(11210) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11210)))) severity failure;
    assert RAM(11211) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11211)))) severity failure;
    assert RAM(11212) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11212)))) severity failure;
    assert RAM(11213) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11213)))) severity failure;
    assert RAM(11214) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11214)))) severity failure;
    assert RAM(11215) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11215)))) severity failure;
    assert RAM(11216) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11216)))) severity failure;
    assert RAM(11217) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11217)))) severity failure;
    assert RAM(11218) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11218)))) severity failure;
    assert RAM(11219) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11219)))) severity failure;
    assert RAM(11220) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11220)))) severity failure;
    assert RAM(11221) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11221)))) severity failure;
    assert RAM(11222) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11222)))) severity failure;
    assert RAM(11223) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11223)))) severity failure;
    assert RAM(11224) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11224)))) severity failure;
    assert RAM(11225) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11225)))) severity failure;
    assert RAM(11226) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11226)))) severity failure;
    assert RAM(11227) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11227)))) severity failure;
    assert RAM(11228) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11228)))) severity failure;
    assert RAM(11229) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11229)))) severity failure;
    assert RAM(11230) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11230)))) severity failure;
    assert RAM(11231) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11231)))) severity failure;
    assert RAM(11232) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11232)))) severity failure;
    assert RAM(11233) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11233)))) severity failure;
    assert RAM(11234) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11234)))) severity failure;
    assert RAM(11235) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11235)))) severity failure;
    assert RAM(11236) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11236)))) severity failure;
    assert RAM(11237) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11237)))) severity failure;
    assert RAM(11238) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11238)))) severity failure;
    assert RAM(11239) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11239)))) severity failure;
    assert RAM(11240) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11240)))) severity failure;
    assert RAM(11241) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11241)))) severity failure;
    assert RAM(11242) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11242)))) severity failure;
    assert RAM(11243) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11243)))) severity failure;
    assert RAM(11244) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11244)))) severity failure;
    assert RAM(11245) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11245)))) severity failure;
    assert RAM(11246) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11246)))) severity failure;
    assert RAM(11247) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11247)))) severity failure;
    assert RAM(11248) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11248)))) severity failure;
    assert RAM(11249) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11249)))) severity failure;
    assert RAM(11250) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11250)))) severity failure;
    assert RAM(11251) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11251)))) severity failure;
    assert RAM(11252) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11252)))) severity failure;
    assert RAM(11253) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11253)))) severity failure;
    assert RAM(11254) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11254)))) severity failure;
    assert RAM(11255) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11255)))) severity failure;
    assert RAM(11256) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11256)))) severity failure;
    assert RAM(11257) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11257)))) severity failure;
    assert RAM(11258) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11258)))) severity failure;
    assert RAM(11259) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11259)))) severity failure;
    assert RAM(11260) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11260)))) severity failure;
    assert RAM(11261) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11261)))) severity failure;
    assert RAM(11262) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11262)))) severity failure;
    assert RAM(11263) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11263)))) severity failure;
    assert RAM(11264) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11264)))) severity failure;
    assert RAM(11265) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11265)))) severity failure;
    assert RAM(11266) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11266)))) severity failure;
    assert RAM(11267) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11267)))) severity failure;
    assert RAM(11268) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11268)))) severity failure;
    assert RAM(11269) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11269)))) severity failure;
    assert RAM(11270) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11270)))) severity failure;
    assert RAM(11271) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11271)))) severity failure;
    assert RAM(11272) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11272)))) severity failure;
    assert RAM(11273) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11273)))) severity failure;
    assert RAM(11274) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11274)))) severity failure;
    assert RAM(11275) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11275)))) severity failure;
    assert RAM(11276) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11276)))) severity failure;
    assert RAM(11277) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11277)))) severity failure;
    assert RAM(11278) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11278)))) severity failure;
    assert RAM(11279) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11279)))) severity failure;
    assert RAM(11280) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11280)))) severity failure;
    assert RAM(11281) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11281)))) severity failure;
    assert RAM(11282) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11282)))) severity failure;
    assert RAM(11283) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11283)))) severity failure;
    assert RAM(11284) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11284)))) severity failure;
    assert RAM(11285) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11285)))) severity failure;
    assert RAM(11286) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11286)))) severity failure;
    assert RAM(11287) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11287)))) severity failure;
    assert RAM(11288) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11288)))) severity failure;
    assert RAM(11289) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11289)))) severity failure;
    assert RAM(11290) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11290)))) severity failure;
    assert RAM(11291) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11291)))) severity failure;
    assert RAM(11292) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11292)))) severity failure;
    assert RAM(11293) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11293)))) severity failure;
    assert RAM(11294) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11294)))) severity failure;
    assert RAM(11295) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11295)))) severity failure;
    assert RAM(11296) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11296)))) severity failure;
    assert RAM(11297) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11297)))) severity failure;
    assert RAM(11298) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11298)))) severity failure;
    assert RAM(11299) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11299)))) severity failure;
    assert RAM(11300) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11300)))) severity failure;
    assert RAM(11301) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11301)))) severity failure;
    assert RAM(11302) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11302)))) severity failure;
    assert RAM(11303) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11303)))) severity failure;
    assert RAM(11304) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11304)))) severity failure;
    assert RAM(11305) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11305)))) severity failure;
    assert RAM(11306) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11306)))) severity failure;
    assert RAM(11307) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11307)))) severity failure;
    assert RAM(11308) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11308)))) severity failure;
    assert RAM(11309) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11309)))) severity failure;
    assert RAM(11310) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11310)))) severity failure;
    assert RAM(11311) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11311)))) severity failure;
    assert RAM(11312) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11312)))) severity failure;
    assert RAM(11313) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11313)))) severity failure;
    assert RAM(11314) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11314)))) severity failure;
    assert RAM(11315) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11315)))) severity failure;
    assert RAM(11316) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11316)))) severity failure;
    assert RAM(11317) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11317)))) severity failure;
    assert RAM(11318) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11318)))) severity failure;
    assert RAM(11319) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11319)))) severity failure;
    assert RAM(11320) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11320)))) severity failure;
    assert RAM(11321) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11321)))) severity failure;
    assert RAM(11322) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11322)))) severity failure;
    assert RAM(11323) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11323)))) severity failure;
    assert RAM(11324) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11324)))) severity failure;
    assert RAM(11325) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11325)))) severity failure;
    assert RAM(11326) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11326)))) severity failure;
    assert RAM(11327) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11327)))) severity failure;
    assert RAM(11328) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11328)))) severity failure;
    assert RAM(11329) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11329)))) severity failure;
    assert RAM(11330) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11330)))) severity failure;
    assert RAM(11331) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11331)))) severity failure;
    assert RAM(11332) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11332)))) severity failure;
    assert RAM(11333) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11333)))) severity failure;
    assert RAM(11334) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11334)))) severity failure;
    assert RAM(11335) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11335)))) severity failure;
    assert RAM(11336) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11336)))) severity failure;
    assert RAM(11337) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11337)))) severity failure;
    assert RAM(11338) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11338)))) severity failure;
    assert RAM(11339) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11339)))) severity failure;
    assert RAM(11340) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11340)))) severity failure;
    assert RAM(11341) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11341)))) severity failure;
    assert RAM(11342) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11342)))) severity failure;
    assert RAM(11343) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11343)))) severity failure;
    assert RAM(11344) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11344)))) severity failure;
    assert RAM(11345) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11345)))) severity failure;
    assert RAM(11346) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11346)))) severity failure;
    assert RAM(11347) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11347)))) severity failure;
    assert RAM(11348) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11348)))) severity failure;
    assert RAM(11349) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11349)))) severity failure;
    assert RAM(11350) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11350)))) severity failure;
    assert RAM(11351) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11351)))) severity failure;
    assert RAM(11352) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11352)))) severity failure;
    assert RAM(11353) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11353)))) severity failure;
    assert RAM(11354) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11354)))) severity failure;
    assert RAM(11355) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11355)))) severity failure;
    assert RAM(11356) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11356)))) severity failure;
    assert RAM(11357) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11357)))) severity failure;
    assert RAM(11358) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11358)))) severity failure;
    assert RAM(11359) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11359)))) severity failure;
    assert RAM(11360) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11360)))) severity failure;
    assert RAM(11361) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11361)))) severity failure;
    assert RAM(11362) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11362)))) severity failure;
    assert RAM(11363) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11363)))) severity failure;
    assert RAM(11364) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11364)))) severity failure;
    assert RAM(11365) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11365)))) severity failure;
    assert RAM(11366) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11366)))) severity failure;
    assert RAM(11367) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11367)))) severity failure;
    assert RAM(11368) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11368)))) severity failure;
    assert RAM(11369) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11369)))) severity failure;
    assert RAM(11370) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11370)))) severity failure;
    assert RAM(11371) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11371)))) severity failure;
    assert RAM(11372) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11372)))) severity failure;
    assert RAM(11373) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11373)))) severity failure;
    assert RAM(11374) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11374)))) severity failure;
    assert RAM(11375) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11375)))) severity failure;
    assert RAM(11376) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11376)))) severity failure;
    assert RAM(11377) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11377)))) severity failure;
    assert RAM(11378) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11378)))) severity failure;
    assert RAM(11379) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11379)))) severity failure;
    assert RAM(11380) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11380)))) severity failure;
    assert RAM(11381) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11381)))) severity failure;
    assert RAM(11382) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11382)))) severity failure;
    assert RAM(11383) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11383)))) severity failure;
    assert RAM(11384) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11384)))) severity failure;
    assert RAM(11385) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11385)))) severity failure;
    assert RAM(11386) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11386)))) severity failure;
    assert RAM(11387) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11387)))) severity failure;
    assert RAM(11388) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11388)))) severity failure;
    assert RAM(11389) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11389)))) severity failure;
    assert RAM(11390) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11390)))) severity failure;
    assert RAM(11391) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11391)))) severity failure;
    assert RAM(11392) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11392)))) severity failure;
    assert RAM(11393) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11393)))) severity failure;
    assert RAM(11394) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11394)))) severity failure;
    assert RAM(11395) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11395)))) severity failure;
    assert RAM(11396) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11396)))) severity failure;
    assert RAM(11397) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11397)))) severity failure;
    assert RAM(11398) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11398)))) severity failure;
    assert RAM(11399) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11399)))) severity failure;
    assert RAM(11400) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11400)))) severity failure;
    assert RAM(11401) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11401)))) severity failure;
    assert RAM(11402) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11402)))) severity failure;
    assert RAM(11403) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11403)))) severity failure;
    assert RAM(11404) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11404)))) severity failure;
    assert RAM(11405) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11405)))) severity failure;
    assert RAM(11406) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11406)))) severity failure;
    assert RAM(11407) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11407)))) severity failure;
    assert RAM(11408) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11408)))) severity failure;
    assert RAM(11409) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11409)))) severity failure;
    assert RAM(11410) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11410)))) severity failure;
    assert RAM(11411) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11411)))) severity failure;
    assert RAM(11412) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11412)))) severity failure;
    assert RAM(11413) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11413)))) severity failure;
    assert RAM(11414) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11414)))) severity failure;
    assert RAM(11415) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11415)))) severity failure;
    assert RAM(11416) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11416)))) severity failure;
    assert RAM(11417) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11417)))) severity failure;
    assert RAM(11418) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11418)))) severity failure;
    assert RAM(11419) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11419)))) severity failure;
    assert RAM(11420) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11420)))) severity failure;
    assert RAM(11421) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11421)))) severity failure;
    assert RAM(11422) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11422)))) severity failure;
    assert RAM(11423) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11423)))) severity failure;
    assert RAM(11424) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11424)))) severity failure;
    assert RAM(11425) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11425)))) severity failure;
    assert RAM(11426) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11426)))) severity failure;
    assert RAM(11427) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11427)))) severity failure;
    assert RAM(11428) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11428)))) severity failure;
    assert RAM(11429) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11429)))) severity failure;
    assert RAM(11430) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11430)))) severity failure;
    assert RAM(11431) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11431)))) severity failure;
    assert RAM(11432) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11432)))) severity failure;
    assert RAM(11433) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11433)))) severity failure;
    assert RAM(11434) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11434)))) severity failure;
    assert RAM(11435) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11435)))) severity failure;
    assert RAM(11436) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11436)))) severity failure;
    assert RAM(11437) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11437)))) severity failure;
    assert RAM(11438) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11438)))) severity failure;
    assert RAM(11439) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11439)))) severity failure;
    assert RAM(11440) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11440)))) severity failure;
    assert RAM(11441) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11441)))) severity failure;
    assert RAM(11442) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11442)))) severity failure;
    assert RAM(11443) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11443)))) severity failure;
    assert RAM(11444) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11444)))) severity failure;
    assert RAM(11445) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11445)))) severity failure;
    assert RAM(11446) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11446)))) severity failure;
    assert RAM(11447) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11447)))) severity failure;
    assert RAM(11448) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11448)))) severity failure;
    assert RAM(11449) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11449)))) severity failure;
    assert RAM(11450) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11450)))) severity failure;
    assert RAM(11451) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11451)))) severity failure;
    assert RAM(11452) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11452)))) severity failure;
    assert RAM(11453) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11453)))) severity failure;
    assert RAM(11454) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11454)))) severity failure;
    assert RAM(11455) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11455)))) severity failure;
    assert RAM(11456) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11456)))) severity failure;
    assert RAM(11457) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11457)))) severity failure;
    assert RAM(11458) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11458)))) severity failure;
    assert RAM(11459) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11459)))) severity failure;
    assert RAM(11460) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11460)))) severity failure;
    assert RAM(11461) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11461)))) severity failure;
    assert RAM(11462) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11462)))) severity failure;
    assert RAM(11463) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11463)))) severity failure;
    assert RAM(11464) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11464)))) severity failure;
    assert RAM(11465) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11465)))) severity failure;
    assert RAM(11466) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11466)))) severity failure;
    assert RAM(11467) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11467)))) severity failure;
    assert RAM(11468) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11468)))) severity failure;
    assert RAM(11469) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11469)))) severity failure;
    assert RAM(11470) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11470)))) severity failure;
    assert RAM(11471) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11471)))) severity failure;
    assert RAM(11472) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11472)))) severity failure;
    assert RAM(11473) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11473)))) severity failure;
    assert RAM(11474) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11474)))) severity failure;
    assert RAM(11475) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11475)))) severity failure;
    assert RAM(11476) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11476)))) severity failure;
    assert RAM(11477) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11477)))) severity failure;
    assert RAM(11478) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11478)))) severity failure;
    assert RAM(11479) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11479)))) severity failure;
    assert RAM(11480) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11480)))) severity failure;
    assert RAM(11481) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11481)))) severity failure;
    assert RAM(11482) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11482)))) severity failure;
    assert RAM(11483) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11483)))) severity failure;
    assert RAM(11484) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11484)))) severity failure;
    assert RAM(11485) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11485)))) severity failure;
    assert RAM(11486) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11486)))) severity failure;
    assert RAM(11487) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11487)))) severity failure;
    assert RAM(11488) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11488)))) severity failure;
    assert RAM(11489) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11489)))) severity failure;
    assert RAM(11490) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11490)))) severity failure;
    assert RAM(11491) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11491)))) severity failure;
    assert RAM(11492) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11492)))) severity failure;
    assert RAM(11493) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11493)))) severity failure;
    assert RAM(11494) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11494)))) severity failure;
    assert RAM(11495) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11495)))) severity failure;
    assert RAM(11496) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11496)))) severity failure;
    assert RAM(11497) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11497)))) severity failure;
    assert RAM(11498) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11498)))) severity failure;
    assert RAM(11499) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11499)))) severity failure;
    assert RAM(11500) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11500)))) severity failure;
    assert RAM(11501) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11501)))) severity failure;
    assert RAM(11502) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11502)))) severity failure;
    assert RAM(11503) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11503)))) severity failure;
    assert RAM(11504) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11504)))) severity failure;
    assert RAM(11505) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11505)))) severity failure;
    assert RAM(11506) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11506)))) severity failure;
    assert RAM(11507) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11507)))) severity failure;
    assert RAM(11508) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11508)))) severity failure;
    assert RAM(11509) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11509)))) severity failure;
    assert RAM(11510) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11510)))) severity failure;
    assert RAM(11511) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11511)))) severity failure;
    assert RAM(11512) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11512)))) severity failure;
    assert RAM(11513) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11513)))) severity failure;
    assert RAM(11514) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11514)))) severity failure;
    assert RAM(11515) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11515)))) severity failure;
    assert RAM(11516) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11516)))) severity failure;
    assert RAM(11517) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11517)))) severity failure;
    assert RAM(11518) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11518)))) severity failure;
    assert RAM(11519) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11519)))) severity failure;
    assert RAM(11520) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11520)))) severity failure;
    assert RAM(11521) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11521)))) severity failure;
    assert RAM(11522) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11522)))) severity failure;
    assert RAM(11523) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11523)))) severity failure;
    assert RAM(11524) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11524)))) severity failure;
    assert RAM(11525) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11525)))) severity failure;
    assert RAM(11526) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11526)))) severity failure;
    assert RAM(11527) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11527)))) severity failure;
    assert RAM(11528) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11528)))) severity failure;
    assert RAM(11529) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11529)))) severity failure;
    assert RAM(11530) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11530)))) severity failure;
    assert RAM(11531) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11531)))) severity failure;
    assert RAM(11532) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11532)))) severity failure;
    assert RAM(11533) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11533)))) severity failure;
    assert RAM(11534) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11534)))) severity failure;
    assert RAM(11535) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11535)))) severity failure;
    assert RAM(11536) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11536)))) severity failure;
    assert RAM(11537) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11537)))) severity failure;
    assert RAM(11538) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11538)))) severity failure;
    assert RAM(11539) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11539)))) severity failure;
    assert RAM(11540) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11540)))) severity failure;
    assert RAM(11541) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11541)))) severity failure;
    assert RAM(11542) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11542)))) severity failure;
    assert RAM(11543) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11543)))) severity failure;
    assert RAM(11544) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11544)))) severity failure;
    assert RAM(11545) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11545)))) severity failure;
    assert RAM(11546) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11546)))) severity failure;
    assert RAM(11547) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11547)))) severity failure;
    assert RAM(11548) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11548)))) severity failure;
    assert RAM(11549) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11549)))) severity failure;
    assert RAM(11550) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11550)))) severity failure;
    assert RAM(11551) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11551)))) severity failure;
    assert RAM(11552) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11552)))) severity failure;
    assert RAM(11553) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11553)))) severity failure;
    assert RAM(11554) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11554)))) severity failure;
    assert RAM(11555) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11555)))) severity failure;
    assert RAM(11556) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11556)))) severity failure;
    assert RAM(11557) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11557)))) severity failure;
    assert RAM(11558) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11558)))) severity failure;
    assert RAM(11559) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11559)))) severity failure;
    assert RAM(11560) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11560)))) severity failure;
    assert RAM(11561) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11561)))) severity failure;
    assert RAM(11562) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11562)))) severity failure;
    assert RAM(11563) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11563)))) severity failure;
    assert RAM(11564) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11564)))) severity failure;
    assert RAM(11565) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11565)))) severity failure;
    assert RAM(11566) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11566)))) severity failure;
    assert RAM(11567) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11567)))) severity failure;
    assert RAM(11568) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11568)))) severity failure;
    assert RAM(11569) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11569)))) severity failure;
    assert RAM(11570) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11570)))) severity failure;
    assert RAM(11571) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11571)))) severity failure;
    assert RAM(11572) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11572)))) severity failure;
    assert RAM(11573) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11573)))) severity failure;
    assert RAM(11574) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11574)))) severity failure;
    assert RAM(11575) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11575)))) severity failure;
    assert RAM(11576) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11576)))) severity failure;
    assert RAM(11577) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11577)))) severity failure;
    assert RAM(11578) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11578)))) severity failure;
    assert RAM(11579) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11579)))) severity failure;
    assert RAM(11580) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11580)))) severity failure;
    assert RAM(11581) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11581)))) severity failure;
    assert RAM(11582) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11582)))) severity failure;
    assert RAM(11583) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11583)))) severity failure;
    assert RAM(11584) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11584)))) severity failure;
    assert RAM(11585) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11585)))) severity failure;
    assert RAM(11586) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11586)))) severity failure;
    assert RAM(11587) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11587)))) severity failure;
    assert RAM(11588) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11588)))) severity failure;
    assert RAM(11589) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11589)))) severity failure;
    assert RAM(11590) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11590)))) severity failure;
    assert RAM(11591) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11591)))) severity failure;
    assert RAM(11592) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11592)))) severity failure;
    assert RAM(11593) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11593)))) severity failure;
    assert RAM(11594) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11594)))) severity failure;
    assert RAM(11595) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11595)))) severity failure;
    assert RAM(11596) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11596)))) severity failure;
    assert RAM(11597) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11597)))) severity failure;
    assert RAM(11598) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11598)))) severity failure;
    assert RAM(11599) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11599)))) severity failure;
    assert RAM(11600) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11600)))) severity failure;
    assert RAM(11601) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11601)))) severity failure;
    assert RAM(11602) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11602)))) severity failure;
    assert RAM(11603) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11603)))) severity failure;
    assert RAM(11604) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11604)))) severity failure;
    assert RAM(11605) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11605)))) severity failure;
    assert RAM(11606) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11606)))) severity failure;
    assert RAM(11607) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11607)))) severity failure;
    assert RAM(11608) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11608)))) severity failure;
    assert RAM(11609) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11609)))) severity failure;
    assert RAM(11610) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11610)))) severity failure;
    assert RAM(11611) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11611)))) severity failure;
    assert RAM(11612) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11612)))) severity failure;
    assert RAM(11613) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11613)))) severity failure;
    assert RAM(11614) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11614)))) severity failure;
    assert RAM(11615) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11615)))) severity failure;
    assert RAM(11616) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11616)))) severity failure;
    assert RAM(11617) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11617)))) severity failure;
    assert RAM(11618) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11618)))) severity failure;
    assert RAM(11619) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11619)))) severity failure;
    assert RAM(11620) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11620)))) severity failure;
    assert RAM(11621) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11621)))) severity failure;
    assert RAM(11622) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11622)))) severity failure;
    assert RAM(11623) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11623)))) severity failure;
    assert RAM(11624) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11624)))) severity failure;
    assert RAM(11625) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11625)))) severity failure;
    assert RAM(11626) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11626)))) severity failure;
    assert RAM(11627) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11627)))) severity failure;
    assert RAM(11628) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11628)))) severity failure;
    assert RAM(11629) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11629)))) severity failure;
    assert RAM(11630) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11630)))) severity failure;
    assert RAM(11631) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11631)))) severity failure;
    assert RAM(11632) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11632)))) severity failure;
    assert RAM(11633) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11633)))) severity failure;
    assert RAM(11634) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11634)))) severity failure;
    assert RAM(11635) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11635)))) severity failure;
    assert RAM(11636) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11636)))) severity failure;
    assert RAM(11637) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11637)))) severity failure;
    assert RAM(11638) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11638)))) severity failure;
    assert RAM(11639) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11639)))) severity failure;
    assert RAM(11640) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11640)))) severity failure;
    assert RAM(11641) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11641)))) severity failure;
    assert RAM(11642) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11642)))) severity failure;
    assert RAM(11643) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11643)))) severity failure;
    assert RAM(11644) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11644)))) severity failure;
    assert RAM(11645) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11645)))) severity failure;
    assert RAM(11646) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11646)))) severity failure;
    assert RAM(11647) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11647)))) severity failure;
    assert RAM(11648) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11648)))) severity failure;
    assert RAM(11649) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11649)))) severity failure;
    assert RAM(11650) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11650)))) severity failure;
    assert RAM(11651) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11651)))) severity failure;
    assert RAM(11652) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11652)))) severity failure;
    assert RAM(11653) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11653)))) severity failure;
    assert RAM(11654) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11654)))) severity failure;
    assert RAM(11655) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11655)))) severity failure;
    assert RAM(11656) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11656)))) severity failure;
    assert RAM(11657) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11657)))) severity failure;
    assert RAM(11658) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11658)))) severity failure;
    assert RAM(11659) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11659)))) severity failure;
    assert RAM(11660) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11660)))) severity failure;
    assert RAM(11661) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11661)))) severity failure;
    assert RAM(11662) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11662)))) severity failure;
    assert RAM(11663) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11663)))) severity failure;
    assert RAM(11664) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11664)))) severity failure;
    assert RAM(11665) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11665)))) severity failure;
    assert RAM(11666) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11666)))) severity failure;
    assert RAM(11667) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11667)))) severity failure;
    assert RAM(11668) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11668)))) severity failure;
    assert RAM(11669) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11669)))) severity failure;
    assert RAM(11670) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11670)))) severity failure;
    assert RAM(11671) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11671)))) severity failure;
    assert RAM(11672) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11672)))) severity failure;
    assert RAM(11673) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11673)))) severity failure;
    assert RAM(11674) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11674)))) severity failure;
    assert RAM(11675) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11675)))) severity failure;
    assert RAM(11676) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11676)))) severity failure;
    assert RAM(11677) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11677)))) severity failure;
    assert RAM(11678) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11678)))) severity failure;
    assert RAM(11679) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11679)))) severity failure;
    assert RAM(11680) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11680)))) severity failure;
    assert RAM(11681) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11681)))) severity failure;
    assert RAM(11682) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11682)))) severity failure;
    assert RAM(11683) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11683)))) severity failure;
    assert RAM(11684) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11684)))) severity failure;
    assert RAM(11685) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11685)))) severity failure;
    assert RAM(11686) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11686)))) severity failure;
    assert RAM(11687) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11687)))) severity failure;
    assert RAM(11688) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11688)))) severity failure;
    assert RAM(11689) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11689)))) severity failure;
    assert RAM(11690) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11690)))) severity failure;
    assert RAM(11691) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11691)))) severity failure;
    assert RAM(11692) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11692)))) severity failure;
    assert RAM(11693) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11693)))) severity failure;
    assert RAM(11694) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11694)))) severity failure;
    assert RAM(11695) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11695)))) severity failure;
    assert RAM(11696) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11696)))) severity failure;
    assert RAM(11697) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11697)))) severity failure;
    assert RAM(11698) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11698)))) severity failure;
    assert RAM(11699) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11699)))) severity failure;
    assert RAM(11700) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11700)))) severity failure;
    assert RAM(11701) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11701)))) severity failure;
    assert RAM(11702) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11702)))) severity failure;
    assert RAM(11703) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11703)))) severity failure;
    assert RAM(11704) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11704)))) severity failure;
    assert RAM(11705) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11705)))) severity failure;
    assert RAM(11706) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11706)))) severity failure;
    assert RAM(11707) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11707)))) severity failure;
    assert RAM(11708) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11708)))) severity failure;
    assert RAM(11709) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11709)))) severity failure;
    assert RAM(11710) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11710)))) severity failure;
    assert RAM(11711) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11711)))) severity failure;
    assert RAM(11712) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11712)))) severity failure;
    assert RAM(11713) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11713)))) severity failure;
    assert RAM(11714) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11714)))) severity failure;
    assert RAM(11715) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11715)))) severity failure;
    assert RAM(11716) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11716)))) severity failure;
    assert RAM(11717) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11717)))) severity failure;
    assert RAM(11718) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11718)))) severity failure;
    assert RAM(11719) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11719)))) severity failure;
    assert RAM(11720) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11720)))) severity failure;
    assert RAM(11721) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11721)))) severity failure;
    assert RAM(11722) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11722)))) severity failure;
    assert RAM(11723) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11723)))) severity failure;
    assert RAM(11724) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11724)))) severity failure;
    assert RAM(11725) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11725)))) severity failure;
    assert RAM(11726) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11726)))) severity failure;
    assert RAM(11727) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11727)))) severity failure;
    assert RAM(11728) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11728)))) severity failure;
    assert RAM(11729) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11729)))) severity failure;
    assert RAM(11730) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11730)))) severity failure;
    assert RAM(11731) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11731)))) severity failure;
    assert RAM(11732) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11732)))) severity failure;
    assert RAM(11733) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11733)))) severity failure;
    assert RAM(11734) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11734)))) severity failure;
    assert RAM(11735) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11735)))) severity failure;
    assert RAM(11736) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11736)))) severity failure;
    assert RAM(11737) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11737)))) severity failure;
    assert RAM(11738) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11738)))) severity failure;
    assert RAM(11739) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11739)))) severity failure;
    assert RAM(11740) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11740)))) severity failure;
    assert RAM(11741) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11741)))) severity failure;
    assert RAM(11742) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11742)))) severity failure;
    assert RAM(11743) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11743)))) severity failure;
    assert RAM(11744) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11744)))) severity failure;
    assert RAM(11745) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11745)))) severity failure;
    assert RAM(11746) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11746)))) severity failure;
    assert RAM(11747) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11747)))) severity failure;
    assert RAM(11748) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11748)))) severity failure;
    assert RAM(11749) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11749)))) severity failure;
    assert RAM(11750) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11750)))) severity failure;
    assert RAM(11751) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11751)))) severity failure;
    assert RAM(11752) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11752)))) severity failure;
    assert RAM(11753) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11753)))) severity failure;
    assert RAM(11754) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11754)))) severity failure;
    assert RAM(11755) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11755)))) severity failure;
    assert RAM(11756) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11756)))) severity failure;
    assert RAM(11757) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11757)))) severity failure;
    assert RAM(11758) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11758)))) severity failure;
    assert RAM(11759) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11759)))) severity failure;
    assert RAM(11760) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11760)))) severity failure;
    assert RAM(11761) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11761)))) severity failure;
    assert RAM(11762) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11762)))) severity failure;
    assert RAM(11763) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11763)))) severity failure;
    assert RAM(11764) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11764)))) severity failure;
    assert RAM(11765) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11765)))) severity failure;
    assert RAM(11766) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11766)))) severity failure;
    assert RAM(11767) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11767)))) severity failure;
    assert RAM(11768) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11768)))) severity failure;
    assert RAM(11769) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11769)))) severity failure;
    assert RAM(11770) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11770)))) severity failure;
    assert RAM(11771) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11771)))) severity failure;
    assert RAM(11772) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11772)))) severity failure;
    assert RAM(11773) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11773)))) severity failure;
    assert RAM(11774) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11774)))) severity failure;
    assert RAM(11775) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11775)))) severity failure;
    assert RAM(11776) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11776)))) severity failure;
    assert RAM(11777) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11777)))) severity failure;
    assert RAM(11778) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11778)))) severity failure;
    assert RAM(11779) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11779)))) severity failure;
    assert RAM(11780) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11780)))) severity failure;
    assert RAM(11781) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11781)))) severity failure;
    assert RAM(11782) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11782)))) severity failure;
    assert RAM(11783) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11783)))) severity failure;
    assert RAM(11784) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11784)))) severity failure;
    assert RAM(11785) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11785)))) severity failure;
    assert RAM(11786) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11786)))) severity failure;
    assert RAM(11787) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11787)))) severity failure;
    assert RAM(11788) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11788)))) severity failure;
    assert RAM(11789) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11789)))) severity failure;
    assert RAM(11790) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11790)))) severity failure;
    assert RAM(11791) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11791)))) severity failure;
    assert RAM(11792) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11792)))) severity failure;
    assert RAM(11793) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11793)))) severity failure;
    assert RAM(11794) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11794)))) severity failure;
    assert RAM(11795) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11795)))) severity failure;
    assert RAM(11796) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11796)))) severity failure;
    assert RAM(11797) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11797)))) severity failure;
    assert RAM(11798) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11798)))) severity failure;
    assert RAM(11799) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11799)))) severity failure;
    assert RAM(11800) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11800)))) severity failure;
    assert RAM(11801) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11801)))) severity failure;
    assert RAM(11802) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11802)))) severity failure;
    assert RAM(11803) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11803)))) severity failure;
    assert RAM(11804) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11804)))) severity failure;
    assert RAM(11805) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11805)))) severity failure;
    assert RAM(11806) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11806)))) severity failure;
    assert RAM(11807) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11807)))) severity failure;
    assert RAM(11808) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11808)))) severity failure;
    assert RAM(11809) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11809)))) severity failure;
    assert RAM(11810) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11810)))) severity failure;
    assert RAM(11811) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11811)))) severity failure;
    assert RAM(11812) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11812)))) severity failure;
    assert RAM(11813) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11813)))) severity failure;
    assert RAM(11814) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11814)))) severity failure;
    assert RAM(11815) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11815)))) severity failure;
    assert RAM(11816) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11816)))) severity failure;
    assert RAM(11817) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11817)))) severity failure;
    assert RAM(11818) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11818)))) severity failure;
    assert RAM(11819) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11819)))) severity failure;
    assert RAM(11820) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11820)))) severity failure;
    assert RAM(11821) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11821)))) severity failure;
    assert RAM(11822) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11822)))) severity failure;
    assert RAM(11823) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11823)))) severity failure;
    assert RAM(11824) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11824)))) severity failure;
    assert RAM(11825) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11825)))) severity failure;
    assert RAM(11826) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11826)))) severity failure;
    assert RAM(11827) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11827)))) severity failure;
    assert RAM(11828) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11828)))) severity failure;
    assert RAM(11829) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11829)))) severity failure;
    assert RAM(11830) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11830)))) severity failure;
    assert RAM(11831) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11831)))) severity failure;
    assert RAM(11832) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11832)))) severity failure;
    assert RAM(11833) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11833)))) severity failure;
    assert RAM(11834) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11834)))) severity failure;
    assert RAM(11835) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11835)))) severity failure;
    assert RAM(11836) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11836)))) severity failure;
    assert RAM(11837) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11837)))) severity failure;
    assert RAM(11838) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11838)))) severity failure;
    assert RAM(11839) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11839)))) severity failure;
    assert RAM(11840) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11840)))) severity failure;
    assert RAM(11841) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11841)))) severity failure;
    assert RAM(11842) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11842)))) severity failure;
    assert RAM(11843) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11843)))) severity failure;
    assert RAM(11844) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11844)))) severity failure;
    assert RAM(11845) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11845)))) severity failure;
    assert RAM(11846) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11846)))) severity failure;
    assert RAM(11847) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11847)))) severity failure;
    assert RAM(11848) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11848)))) severity failure;
    assert RAM(11849) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11849)))) severity failure;
    assert RAM(11850) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11850)))) severity failure;
    assert RAM(11851) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11851)))) severity failure;
    assert RAM(11852) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11852)))) severity failure;
    assert RAM(11853) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11853)))) severity failure;
    assert RAM(11854) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11854)))) severity failure;
    assert RAM(11855) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11855)))) severity failure;
    assert RAM(11856) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11856)))) severity failure;
    assert RAM(11857) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11857)))) severity failure;
    assert RAM(11858) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11858)))) severity failure;
    assert RAM(11859) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11859)))) severity failure;
    assert RAM(11860) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11860)))) severity failure;
    assert RAM(11861) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11861)))) severity failure;
    assert RAM(11862) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11862)))) severity failure;
    assert RAM(11863) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11863)))) severity failure;
    assert RAM(11864) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11864)))) severity failure;
    assert RAM(11865) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11865)))) severity failure;
    assert RAM(11866) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11866)))) severity failure;
    assert RAM(11867) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11867)))) severity failure;
    assert RAM(11868) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11868)))) severity failure;
    assert RAM(11869) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11869)))) severity failure;
    assert RAM(11870) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11870)))) severity failure;
    assert RAM(11871) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11871)))) severity failure;
    assert RAM(11872) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11872)))) severity failure;
    assert RAM(11873) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11873)))) severity failure;
    assert RAM(11874) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11874)))) severity failure;
    assert RAM(11875) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11875)))) severity failure;
    assert RAM(11876) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11876)))) severity failure;
    assert RAM(11877) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11877)))) severity failure;
    assert RAM(11878) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11878)))) severity failure;
    assert RAM(11879) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11879)))) severity failure;
    assert RAM(11880) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11880)))) severity failure;
    assert RAM(11881) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11881)))) severity failure;
    assert RAM(11882) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11882)))) severity failure;
    assert RAM(11883) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11883)))) severity failure;
    assert RAM(11884) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11884)))) severity failure;
    assert RAM(11885) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11885)))) severity failure;
    assert RAM(11886) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11886)))) severity failure;
    assert RAM(11887) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11887)))) severity failure;
    assert RAM(11888) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11888)))) severity failure;
    assert RAM(11889) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11889)))) severity failure;
    assert RAM(11890) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11890)))) severity failure;
    assert RAM(11891) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11891)))) severity failure;
    assert RAM(11892) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11892)))) severity failure;
    assert RAM(11893) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11893)))) severity failure;
    assert RAM(11894) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11894)))) severity failure;
    assert RAM(11895) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11895)))) severity failure;
    assert RAM(11896) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11896)))) severity failure;
    assert RAM(11897) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11897)))) severity failure;
    assert RAM(11898) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11898)))) severity failure;
    assert RAM(11899) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11899)))) severity failure;
    assert RAM(11900) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11900)))) severity failure;
    assert RAM(11901) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11901)))) severity failure;
    assert RAM(11902) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11902)))) severity failure;
    assert RAM(11903) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11903)))) severity failure;
    assert RAM(11904) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11904)))) severity failure;
    assert RAM(11905) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11905)))) severity failure;
    assert RAM(11906) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11906)))) severity failure;
    assert RAM(11907) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11907)))) severity failure;
    assert RAM(11908) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11908)))) severity failure;
    assert RAM(11909) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11909)))) severity failure;
    assert RAM(11910) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11910)))) severity failure;
    assert RAM(11911) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11911)))) severity failure;
    assert RAM(11912) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11912)))) severity failure;
    assert RAM(11913) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11913)))) severity failure;
    assert RAM(11914) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11914)))) severity failure;
    assert RAM(11915) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11915)))) severity failure;
    assert RAM(11916) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11916)))) severity failure;
    assert RAM(11917) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11917)))) severity failure;
    assert RAM(11918) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11918)))) severity failure;
    assert RAM(11919) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11919)))) severity failure;
    assert RAM(11920) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11920)))) severity failure;
    assert RAM(11921) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11921)))) severity failure;
    assert RAM(11922) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11922)))) severity failure;
    assert RAM(11923) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11923)))) severity failure;
    assert RAM(11924) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11924)))) severity failure;
    assert RAM(11925) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11925)))) severity failure;
    assert RAM(11926) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11926)))) severity failure;
    assert RAM(11927) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11927)))) severity failure;
    assert RAM(11928) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11928)))) severity failure;
    assert RAM(11929) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11929)))) severity failure;
    assert RAM(11930) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11930)))) severity failure;
    assert RAM(11931) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11931)))) severity failure;
    assert RAM(11932) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11932)))) severity failure;
    assert RAM(11933) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11933)))) severity failure;
    assert RAM(11934) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11934)))) severity failure;
    assert RAM(11935) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11935)))) severity failure;
    assert RAM(11936) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11936)))) severity failure;
    assert RAM(11937) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11937)))) severity failure;
    assert RAM(11938) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11938)))) severity failure;
    assert RAM(11939) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11939)))) severity failure;
    assert RAM(11940) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11940)))) severity failure;
    assert RAM(11941) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11941)))) severity failure;
    assert RAM(11942) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11942)))) severity failure;
    assert RAM(11943) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11943)))) severity failure;
    assert RAM(11944) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11944)))) severity failure;
    assert RAM(11945) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11945)))) severity failure;
    assert RAM(11946) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11946)))) severity failure;
    assert RAM(11947) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11947)))) severity failure;
    assert RAM(11948) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11948)))) severity failure;
    assert RAM(11949) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11949)))) severity failure;
    assert RAM(11950) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11950)))) severity failure;
    assert RAM(11951) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11951)))) severity failure;
    assert RAM(11952) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11952)))) severity failure;
    assert RAM(11953) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11953)))) severity failure;
    assert RAM(11954) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11954)))) severity failure;
    assert RAM(11955) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11955)))) severity failure;
    assert RAM(11956) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11956)))) severity failure;
    assert RAM(11957) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11957)))) severity failure;
    assert RAM(11958) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11958)))) severity failure;
    assert RAM(11959) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11959)))) severity failure;
    assert RAM(11960) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11960)))) severity failure;
    assert RAM(11961) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11961)))) severity failure;
    assert RAM(11962) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11962)))) severity failure;
    assert RAM(11963) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11963)))) severity failure;
    assert RAM(11964) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11964)))) severity failure;
    assert RAM(11965) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11965)))) severity failure;
    assert RAM(11966) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11966)))) severity failure;
    assert RAM(11967) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11967)))) severity failure;
    assert RAM(11968) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11968)))) severity failure;
    assert RAM(11969) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11969)))) severity failure;
    assert RAM(11970) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11970)))) severity failure;
    assert RAM(11971) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11971)))) severity failure;
    assert RAM(11972) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11972)))) severity failure;
    assert RAM(11973) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11973)))) severity failure;
    assert RAM(11974) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11974)))) severity failure;
    assert RAM(11975) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11975)))) severity failure;
    assert RAM(11976) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11976)))) severity failure;
    assert RAM(11977) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11977)))) severity failure;
    assert RAM(11978) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11978)))) severity failure;
    assert RAM(11979) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11979)))) severity failure;
    assert RAM(11980) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11980)))) severity failure;
    assert RAM(11981) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11981)))) severity failure;
    assert RAM(11982) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11982)))) severity failure;
    assert RAM(11983) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11983)))) severity failure;
    assert RAM(11984) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11984)))) severity failure;
    assert RAM(11985) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11985)))) severity failure;
    assert RAM(11986) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11986)))) severity failure;
    assert RAM(11987) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11987)))) severity failure;
    assert RAM(11988) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11988)))) severity failure;
    assert RAM(11989) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11989)))) severity failure;
    assert RAM(11990) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11990)))) severity failure;
    assert RAM(11991) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11991)))) severity failure;
    assert RAM(11992) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11992)))) severity failure;
    assert RAM(11993) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11993)))) severity failure;
    assert RAM(11994) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11994)))) severity failure;
    assert RAM(11995) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11995)))) severity failure;
    assert RAM(11996) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11996)))) severity failure;
    assert RAM(11997) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11997)))) severity failure;
    assert RAM(11998) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(11998)))) severity failure;
    assert RAM(11999) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(11999)))) severity failure;
    assert RAM(12000) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12000)))) severity failure;
    assert RAM(12001) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12001)))) severity failure;
    assert RAM(12002) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12002)))) severity failure;
    assert RAM(12003) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12003)))) severity failure;
    assert RAM(12004) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12004)))) severity failure;
    assert RAM(12005) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12005)))) severity failure;
    assert RAM(12006) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12006)))) severity failure;
    assert RAM(12007) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12007)))) severity failure;
    assert RAM(12008) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12008)))) severity failure;
    assert RAM(12009) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12009)))) severity failure;
    assert RAM(12010) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12010)))) severity failure;
    assert RAM(12011) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12011)))) severity failure;
    assert RAM(12012) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12012)))) severity failure;
    assert RAM(12013) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12013)))) severity failure;
    assert RAM(12014) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12014)))) severity failure;
    assert RAM(12015) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12015)))) severity failure;
    assert RAM(12016) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12016)))) severity failure;
    assert RAM(12017) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12017)))) severity failure;
    assert RAM(12018) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12018)))) severity failure;
    assert RAM(12019) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12019)))) severity failure;
    assert RAM(12020) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12020)))) severity failure;
    assert RAM(12021) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12021)))) severity failure;
    assert RAM(12022) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12022)))) severity failure;
    assert RAM(12023) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12023)))) severity failure;
    assert RAM(12024) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12024)))) severity failure;
    assert RAM(12025) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12025)))) severity failure;
    assert RAM(12026) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12026)))) severity failure;
    assert RAM(12027) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12027)))) severity failure;
    assert RAM(12028) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12028)))) severity failure;
    assert RAM(12029) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12029)))) severity failure;
    assert RAM(12030) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12030)))) severity failure;
    assert RAM(12031) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12031)))) severity failure;
    assert RAM(12032) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12032)))) severity failure;
    assert RAM(12033) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12033)))) severity failure;
    assert RAM(12034) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12034)))) severity failure;
    assert RAM(12035) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12035)))) severity failure;
    assert RAM(12036) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12036)))) severity failure;
    assert RAM(12037) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12037)))) severity failure;
    assert RAM(12038) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12038)))) severity failure;
    assert RAM(12039) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12039)))) severity failure;
    assert RAM(12040) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12040)))) severity failure;
    assert RAM(12041) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12041)))) severity failure;
    assert RAM(12042) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12042)))) severity failure;
    assert RAM(12043) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12043)))) severity failure;
    assert RAM(12044) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12044)))) severity failure;
    assert RAM(12045) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12045)))) severity failure;
    assert RAM(12046) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12046)))) severity failure;
    assert RAM(12047) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12047)))) severity failure;
    assert RAM(12048) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12048)))) severity failure;
    assert RAM(12049) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12049)))) severity failure;
    assert RAM(12050) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12050)))) severity failure;
    assert RAM(12051) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12051)))) severity failure;
    assert RAM(12052) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12052)))) severity failure;
    assert RAM(12053) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12053)))) severity failure;
    assert RAM(12054) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12054)))) severity failure;
    assert RAM(12055) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12055)))) severity failure;
    assert RAM(12056) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12056)))) severity failure;
    assert RAM(12057) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12057)))) severity failure;
    assert RAM(12058) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12058)))) severity failure;
    assert RAM(12059) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12059)))) severity failure;
    assert RAM(12060) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12060)))) severity failure;
    assert RAM(12061) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12061)))) severity failure;
    assert RAM(12062) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12062)))) severity failure;
    assert RAM(12063) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12063)))) severity failure;
    assert RAM(12064) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12064)))) severity failure;
    assert RAM(12065) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12065)))) severity failure;
    assert RAM(12066) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12066)))) severity failure;
    assert RAM(12067) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12067)))) severity failure;
    assert RAM(12068) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12068)))) severity failure;
    assert RAM(12069) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12069)))) severity failure;
    assert RAM(12070) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12070)))) severity failure;
    assert RAM(12071) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12071)))) severity failure;
    assert RAM(12072) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12072)))) severity failure;
    assert RAM(12073) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12073)))) severity failure;
    assert RAM(12074) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12074)))) severity failure;
    assert RAM(12075) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12075)))) severity failure;
    assert RAM(12076) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12076)))) severity failure;
    assert RAM(12077) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12077)))) severity failure;
    assert RAM(12078) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12078)))) severity failure;
    assert RAM(12079) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12079)))) severity failure;
    assert RAM(12080) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12080)))) severity failure;
    assert RAM(12081) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12081)))) severity failure;
    assert RAM(12082) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12082)))) severity failure;
    assert RAM(12083) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12083)))) severity failure;
    assert RAM(12084) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12084)))) severity failure;
    assert RAM(12085) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12085)))) severity failure;
    assert RAM(12086) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12086)))) severity failure;
    assert RAM(12087) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12087)))) severity failure;
    assert RAM(12088) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12088)))) severity failure;
    assert RAM(12089) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12089)))) severity failure;
    assert RAM(12090) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12090)))) severity failure;
    assert RAM(12091) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12091)))) severity failure;
    assert RAM(12092) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12092)))) severity failure;
    assert RAM(12093) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12093)))) severity failure;
    assert RAM(12094) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12094)))) severity failure;
    assert RAM(12095) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12095)))) severity failure;
    assert RAM(12096) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12096)))) severity failure;
    assert RAM(12097) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12097)))) severity failure;
    assert RAM(12098) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12098)))) severity failure;
    assert RAM(12099) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12099)))) severity failure;
    assert RAM(12100) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12100)))) severity failure;
    assert RAM(12101) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12101)))) severity failure;
    assert RAM(12102) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12102)))) severity failure;
    assert RAM(12103) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12103)))) severity failure;
    assert RAM(12104) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12104)))) severity failure;
    assert RAM(12105) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12105)))) severity failure;
    assert RAM(12106) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12106)))) severity failure;
    assert RAM(12107) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12107)))) severity failure;
    assert RAM(12108) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12108)))) severity failure;
    assert RAM(12109) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12109)))) severity failure;
    assert RAM(12110) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12110)))) severity failure;
    assert RAM(12111) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12111)))) severity failure;
    assert RAM(12112) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12112)))) severity failure;
    assert RAM(12113) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12113)))) severity failure;
    assert RAM(12114) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12114)))) severity failure;
    assert RAM(12115) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12115)))) severity failure;
    assert RAM(12116) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12116)))) severity failure;
    assert RAM(12117) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12117)))) severity failure;
    assert RAM(12118) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12118)))) severity failure;
    assert RAM(12119) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12119)))) severity failure;
    assert RAM(12120) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12120)))) severity failure;
    assert RAM(12121) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12121)))) severity failure;
    assert RAM(12122) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12122)))) severity failure;
    assert RAM(12123) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12123)))) severity failure;
    assert RAM(12124) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12124)))) severity failure;
    assert RAM(12125) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12125)))) severity failure;
    assert RAM(12126) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12126)))) severity failure;
    assert RAM(12127) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12127)))) severity failure;
    assert RAM(12128) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12128)))) severity failure;
    assert RAM(12129) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12129)))) severity failure;
    assert RAM(12130) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12130)))) severity failure;
    assert RAM(12131) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12131)))) severity failure;
    assert RAM(12132) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12132)))) severity failure;
    assert RAM(12133) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12133)))) severity failure;
    assert RAM(12134) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12134)))) severity failure;
    assert RAM(12135) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12135)))) severity failure;
    assert RAM(12136) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12136)))) severity failure;
    assert RAM(12137) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12137)))) severity failure;
    assert RAM(12138) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12138)))) severity failure;
    assert RAM(12139) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12139)))) severity failure;
    assert RAM(12140) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12140)))) severity failure;
    assert RAM(12141) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12141)))) severity failure;
    assert RAM(12142) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12142)))) severity failure;
    assert RAM(12143) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12143)))) severity failure;
    assert RAM(12144) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12144)))) severity failure;
    assert RAM(12145) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12145)))) severity failure;
    assert RAM(12146) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12146)))) severity failure;
    assert RAM(12147) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12147)))) severity failure;
    assert RAM(12148) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12148)))) severity failure;
    assert RAM(12149) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12149)))) severity failure;
    assert RAM(12150) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12150)))) severity failure;
    assert RAM(12151) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12151)))) severity failure;
    assert RAM(12152) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12152)))) severity failure;
    assert RAM(12153) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12153)))) severity failure;
    assert RAM(12154) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12154)))) severity failure;
    assert RAM(12155) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12155)))) severity failure;
    assert RAM(12156) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12156)))) severity failure;
    assert RAM(12157) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12157)))) severity failure;
    assert RAM(12158) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12158)))) severity failure;
    assert RAM(12159) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12159)))) severity failure;
    assert RAM(12160) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12160)))) severity failure;
    assert RAM(12161) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12161)))) severity failure;
    assert RAM(12162) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12162)))) severity failure;
    assert RAM(12163) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12163)))) severity failure;
    assert RAM(12164) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12164)))) severity failure;
    assert RAM(12165) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12165)))) severity failure;
    assert RAM(12166) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12166)))) severity failure;
    assert RAM(12167) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12167)))) severity failure;
    assert RAM(12168) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12168)))) severity failure;
    assert RAM(12169) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12169)))) severity failure;
    assert RAM(12170) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12170)))) severity failure;
    assert RAM(12171) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12171)))) severity failure;
    assert RAM(12172) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12172)))) severity failure;
    assert RAM(12173) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12173)))) severity failure;
    assert RAM(12174) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12174)))) severity failure;
    assert RAM(12175) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12175)))) severity failure;
    assert RAM(12176) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12176)))) severity failure;
    assert RAM(12177) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12177)))) severity failure;
    assert RAM(12178) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12178)))) severity failure;
    assert RAM(12179) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12179)))) severity failure;
    assert RAM(12180) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12180)))) severity failure;
    assert RAM(12181) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12181)))) severity failure;
    assert RAM(12182) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12182)))) severity failure;
    assert RAM(12183) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12183)))) severity failure;
    assert RAM(12184) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12184)))) severity failure;
    assert RAM(12185) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12185)))) severity failure;
    assert RAM(12186) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12186)))) severity failure;
    assert RAM(12187) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12187)))) severity failure;
    assert RAM(12188) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12188)))) severity failure;
    assert RAM(12189) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12189)))) severity failure;
    assert RAM(12190) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12190)))) severity failure;
    assert RAM(12191) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12191)))) severity failure;
    assert RAM(12192) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12192)))) severity failure;
    assert RAM(12193) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12193)))) severity failure;
    assert RAM(12194) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12194)))) severity failure;
    assert RAM(12195) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12195)))) severity failure;
    assert RAM(12196) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12196)))) severity failure;
    assert RAM(12197) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12197)))) severity failure;
    assert RAM(12198) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12198)))) severity failure;
    assert RAM(12199) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12199)))) severity failure;
    assert RAM(12200) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12200)))) severity failure;
    assert RAM(12201) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12201)))) severity failure;
    assert RAM(12202) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12202)))) severity failure;
    assert RAM(12203) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12203)))) severity failure;
    assert RAM(12204) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12204)))) severity failure;
    assert RAM(12205) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12205)))) severity failure;
    assert RAM(12206) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12206)))) severity failure;
    assert RAM(12207) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12207)))) severity failure;
    assert RAM(12208) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12208)))) severity failure;
    assert RAM(12209) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12209)))) severity failure;
    assert RAM(12210) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12210)))) severity failure;
    assert RAM(12211) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12211)))) severity failure;
    assert RAM(12212) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12212)))) severity failure;
    assert RAM(12213) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12213)))) severity failure;
    assert RAM(12214) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12214)))) severity failure;
    assert RAM(12215) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12215)))) severity failure;
    assert RAM(12216) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12216)))) severity failure;
    assert RAM(12217) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12217)))) severity failure;
    assert RAM(12218) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12218)))) severity failure;
    assert RAM(12219) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12219)))) severity failure;
    assert RAM(12220) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12220)))) severity failure;
    assert RAM(12221) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12221)))) severity failure;
    assert RAM(12222) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12222)))) severity failure;
    assert RAM(12223) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12223)))) severity failure;
    assert RAM(12224) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12224)))) severity failure;
    assert RAM(12225) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12225)))) severity failure;
    assert RAM(12226) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12226)))) severity failure;
    assert RAM(12227) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12227)))) severity failure;
    assert RAM(12228) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12228)))) severity failure;
    assert RAM(12229) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12229)))) severity failure;
    assert RAM(12230) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12230)))) severity failure;
    assert RAM(12231) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12231)))) severity failure;
    assert RAM(12232) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12232)))) severity failure;
    assert RAM(12233) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12233)))) severity failure;
    assert RAM(12234) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12234)))) severity failure;
    assert RAM(12235) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12235)))) severity failure;
    assert RAM(12236) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12236)))) severity failure;
    assert RAM(12237) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12237)))) severity failure;
    assert RAM(12238) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12238)))) severity failure;
    assert RAM(12239) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12239)))) severity failure;
    assert RAM(12240) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12240)))) severity failure;
    assert RAM(12241) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12241)))) severity failure;
    assert RAM(12242) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12242)))) severity failure;
    assert RAM(12243) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12243)))) severity failure;
    assert RAM(12244) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12244)))) severity failure;
    assert RAM(12245) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12245)))) severity failure;
    assert RAM(12246) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12246)))) severity failure;
    assert RAM(12247) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12247)))) severity failure;
    assert RAM(12248) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12248)))) severity failure;
    assert RAM(12249) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12249)))) severity failure;
    assert RAM(12250) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12250)))) severity failure;
    assert RAM(12251) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12251)))) severity failure;
    assert RAM(12252) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12252)))) severity failure;
    assert RAM(12253) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12253)))) severity failure;
    assert RAM(12254) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12254)))) severity failure;
    assert RAM(12255) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12255)))) severity failure;
    assert RAM(12256) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12256)))) severity failure;
    assert RAM(12257) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12257)))) severity failure;
    assert RAM(12258) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12258)))) severity failure;
    assert RAM(12259) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12259)))) severity failure;
    assert RAM(12260) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12260)))) severity failure;
    assert RAM(12261) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12261)))) severity failure;
    assert RAM(12262) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12262)))) severity failure;
    assert RAM(12263) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12263)))) severity failure;
    assert RAM(12264) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12264)))) severity failure;
    assert RAM(12265) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12265)))) severity failure;
    assert RAM(12266) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12266)))) severity failure;
    assert RAM(12267) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12267)))) severity failure;
    assert RAM(12268) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12268)))) severity failure;
    assert RAM(12269) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12269)))) severity failure;
    assert RAM(12270) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12270)))) severity failure;
    assert RAM(12271) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12271)))) severity failure;
    assert RAM(12272) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12272)))) severity failure;
    assert RAM(12273) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12273)))) severity failure;
    assert RAM(12274) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12274)))) severity failure;
    assert RAM(12275) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12275)))) severity failure;
    assert RAM(12276) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12276)))) severity failure;
    assert RAM(12277) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12277)))) severity failure;
    assert RAM(12278) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12278)))) severity failure;
    assert RAM(12279) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12279)))) severity failure;
    assert RAM(12280) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12280)))) severity failure;
    assert RAM(12281) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12281)))) severity failure;
    assert RAM(12282) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12282)))) severity failure;
    assert RAM(12283) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12283)))) severity failure;
    assert RAM(12284) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12284)))) severity failure;
    assert RAM(12285) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12285)))) severity failure;
    assert RAM(12286) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12286)))) severity failure;
    assert RAM(12287) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12287)))) severity failure;
    assert RAM(12288) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12288)))) severity failure;
    assert RAM(12289) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12289)))) severity failure;
    assert RAM(12290) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12290)))) severity failure;
    assert RAM(12291) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12291)))) severity failure;
    assert RAM(12292) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12292)))) severity failure;
    assert RAM(12293) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12293)))) severity failure;
    assert RAM(12294) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12294)))) severity failure;
    assert RAM(12295) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12295)))) severity failure;
    assert RAM(12296) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12296)))) severity failure;
    assert RAM(12297) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12297)))) severity failure;
    assert RAM(12298) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12298)))) severity failure;
    assert RAM(12299) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12299)))) severity failure;
    assert RAM(12300) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12300)))) severity failure;
    assert RAM(12301) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12301)))) severity failure;
    assert RAM(12302) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12302)))) severity failure;
    assert RAM(12303) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12303)))) severity failure;
    assert RAM(12304) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12304)))) severity failure;
    assert RAM(12305) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12305)))) severity failure;
    assert RAM(12306) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12306)))) severity failure;
    assert RAM(12307) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12307)))) severity failure;
    assert RAM(12308) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12308)))) severity failure;
    assert RAM(12309) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12309)))) severity failure;
    assert RAM(12310) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12310)))) severity failure;
    assert RAM(12311) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12311)))) severity failure;
    assert RAM(12312) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12312)))) severity failure;
    assert RAM(12313) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12313)))) severity failure;
    assert RAM(12314) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12314)))) severity failure;
    assert RAM(12315) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12315)))) severity failure;
    assert RAM(12316) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12316)))) severity failure;
    assert RAM(12317) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12317)))) severity failure;
    assert RAM(12318) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12318)))) severity failure;
    assert RAM(12319) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12319)))) severity failure;
    assert RAM(12320) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12320)))) severity failure;
    assert RAM(12321) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12321)))) severity failure;
    assert RAM(12322) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12322)))) severity failure;
    assert RAM(12323) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12323)))) severity failure;
    assert RAM(12324) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12324)))) severity failure;
    assert RAM(12325) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12325)))) severity failure;
    assert RAM(12326) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12326)))) severity failure;
    assert RAM(12327) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12327)))) severity failure;
    assert RAM(12328) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12328)))) severity failure;
    assert RAM(12329) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12329)))) severity failure;
    assert RAM(12330) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12330)))) severity failure;
    assert RAM(12331) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12331)))) severity failure;
    assert RAM(12332) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12332)))) severity failure;
    assert RAM(12333) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12333)))) severity failure;
    assert RAM(12334) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12334)))) severity failure;
    assert RAM(12335) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12335)))) severity failure;
    assert RAM(12336) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12336)))) severity failure;
    assert RAM(12337) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12337)))) severity failure;
    assert RAM(12338) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12338)))) severity failure;
    assert RAM(12339) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12339)))) severity failure;
    assert RAM(12340) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12340)))) severity failure;
    assert RAM(12341) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12341)))) severity failure;
    assert RAM(12342) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12342)))) severity failure;
    assert RAM(12343) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12343)))) severity failure;
    assert RAM(12344) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12344)))) severity failure;
    assert RAM(12345) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12345)))) severity failure;
    assert RAM(12346) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12346)))) severity failure;
    assert RAM(12347) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12347)))) severity failure;
    assert RAM(12348) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12348)))) severity failure;
    assert RAM(12349) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12349)))) severity failure;
    assert RAM(12350) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12350)))) severity failure;
    assert RAM(12351) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12351)))) severity failure;
    assert RAM(12352) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12352)))) severity failure;
    assert RAM(12353) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12353)))) severity failure;
    assert RAM(12354) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12354)))) severity failure;
    assert RAM(12355) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12355)))) severity failure;
    assert RAM(12356) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12356)))) severity failure;
    assert RAM(12357) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12357)))) severity failure;
    assert RAM(12358) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12358)))) severity failure;
    assert RAM(12359) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12359)))) severity failure;
    assert RAM(12360) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12360)))) severity failure;
    assert RAM(12361) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12361)))) severity failure;
    assert RAM(12362) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12362)))) severity failure;
    assert RAM(12363) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12363)))) severity failure;
    assert RAM(12364) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12364)))) severity failure;
    assert RAM(12365) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12365)))) severity failure;
    assert RAM(12366) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12366)))) severity failure;
    assert RAM(12367) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12367)))) severity failure;
    assert RAM(12368) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12368)))) severity failure;
    assert RAM(12369) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12369)))) severity failure;
    assert RAM(12370) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12370)))) severity failure;
    assert RAM(12371) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12371)))) severity failure;
    assert RAM(12372) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12372)))) severity failure;
    assert RAM(12373) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12373)))) severity failure;
    assert RAM(12374) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12374)))) severity failure;
    assert RAM(12375) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12375)))) severity failure;
    assert RAM(12376) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12376)))) severity failure;
    assert RAM(12377) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12377)))) severity failure;
    assert RAM(12378) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12378)))) severity failure;
    assert RAM(12379) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12379)))) severity failure;
    assert RAM(12380) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12380)))) severity failure;
    assert RAM(12381) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12381)))) severity failure;
    assert RAM(12382) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12382)))) severity failure;
    assert RAM(12383) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12383)))) severity failure;
    assert RAM(12384) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12384)))) severity failure;
    assert RAM(12385) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12385)))) severity failure;
    assert RAM(12386) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12386)))) severity failure;
    assert RAM(12387) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12387)))) severity failure;
    assert RAM(12388) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12388)))) severity failure;
    assert RAM(12389) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12389)))) severity failure;
    assert RAM(12390) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12390)))) severity failure;
    assert RAM(12391) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12391)))) severity failure;
    assert RAM(12392) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12392)))) severity failure;
    assert RAM(12393) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12393)))) severity failure;
    assert RAM(12394) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12394)))) severity failure;
    assert RAM(12395) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12395)))) severity failure;
    assert RAM(12396) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12396)))) severity failure;
    assert RAM(12397) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12397)))) severity failure;
    assert RAM(12398) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12398)))) severity failure;
    assert RAM(12399) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12399)))) severity failure;
    assert RAM(12400) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12400)))) severity failure;
    assert RAM(12401) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12401)))) severity failure;
    assert RAM(12402) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12402)))) severity failure;
    assert RAM(12403) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12403)))) severity failure;
    assert RAM(12404) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12404)))) severity failure;
    assert RAM(12405) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12405)))) severity failure;
    assert RAM(12406) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12406)))) severity failure;
    assert RAM(12407) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12407)))) severity failure;
    assert RAM(12408) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12408)))) severity failure;
    assert RAM(12409) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12409)))) severity failure;
    assert RAM(12410) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12410)))) severity failure;
    assert RAM(12411) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12411)))) severity failure;
    assert RAM(12412) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12412)))) severity failure;
    assert RAM(12413) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12413)))) severity failure;
    assert RAM(12414) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12414)))) severity failure;
    assert RAM(12415) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12415)))) severity failure;
    assert RAM(12416) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12416)))) severity failure;
    assert RAM(12417) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12417)))) severity failure;
    assert RAM(12418) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12418)))) severity failure;
    assert RAM(12419) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12419)))) severity failure;
    assert RAM(12420) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12420)))) severity failure;
    assert RAM(12421) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12421)))) severity failure;
    assert RAM(12422) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12422)))) severity failure;
    assert RAM(12423) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12423)))) severity failure;
    assert RAM(12424) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12424)))) severity failure;
    assert RAM(12425) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12425)))) severity failure;
    assert RAM(12426) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12426)))) severity failure;
    assert RAM(12427) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12427)))) severity failure;
    assert RAM(12428) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12428)))) severity failure;
    assert RAM(12429) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12429)))) severity failure;
    assert RAM(12430) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12430)))) severity failure;
    assert RAM(12431) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12431)))) severity failure;
    assert RAM(12432) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12432)))) severity failure;
    assert RAM(12433) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12433)))) severity failure;
    assert RAM(12434) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12434)))) severity failure;
    assert RAM(12435) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12435)))) severity failure;
    assert RAM(12436) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12436)))) severity failure;
    assert RAM(12437) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12437)))) severity failure;
    assert RAM(12438) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12438)))) severity failure;
    assert RAM(12439) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12439)))) severity failure;
    assert RAM(12440) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12440)))) severity failure;
    assert RAM(12441) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12441)))) severity failure;
    assert RAM(12442) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12442)))) severity failure;
    assert RAM(12443) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12443)))) severity failure;
    assert RAM(12444) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12444)))) severity failure;
    assert RAM(12445) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12445)))) severity failure;
    assert RAM(12446) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12446)))) severity failure;
    assert RAM(12447) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12447)))) severity failure;
    assert RAM(12448) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12448)))) severity failure;
    assert RAM(12449) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12449)))) severity failure;
    assert RAM(12450) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12450)))) severity failure;
    assert RAM(12451) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12451)))) severity failure;
    assert RAM(12452) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12452)))) severity failure;
    assert RAM(12453) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12453)))) severity failure;
    assert RAM(12454) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12454)))) severity failure;
    assert RAM(12455) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12455)))) severity failure;
    assert RAM(12456) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12456)))) severity failure;
    assert RAM(12457) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12457)))) severity failure;
    assert RAM(12458) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12458)))) severity failure;
    assert RAM(12459) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12459)))) severity failure;
    assert RAM(12460) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12460)))) severity failure;
    assert RAM(12461) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12461)))) severity failure;
    assert RAM(12462) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12462)))) severity failure;
    assert RAM(12463) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12463)))) severity failure;
    assert RAM(12464) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12464)))) severity failure;
    assert RAM(12465) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12465)))) severity failure;
    assert RAM(12466) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12466)))) severity failure;
    assert RAM(12467) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12467)))) severity failure;
    assert RAM(12468) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12468)))) severity failure;
    assert RAM(12469) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12469)))) severity failure;
    assert RAM(12470) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12470)))) severity failure;
    assert RAM(12471) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12471)))) severity failure;
    assert RAM(12472) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12472)))) severity failure;
    assert RAM(12473) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12473)))) severity failure;
    assert RAM(12474) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12474)))) severity failure;
    assert RAM(12475) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12475)))) severity failure;
    assert RAM(12476) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12476)))) severity failure;
    assert RAM(12477) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12477)))) severity failure;
    assert RAM(12478) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12478)))) severity failure;
    assert RAM(12479) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12479)))) severity failure;
    assert RAM(12480) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12480)))) severity failure;
    assert RAM(12481) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12481)))) severity failure;
    assert RAM(12482) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12482)))) severity failure;
    assert RAM(12483) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12483)))) severity failure;
    assert RAM(12484) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12484)))) severity failure;
    assert RAM(12485) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12485)))) severity failure;
    assert RAM(12486) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12486)))) severity failure;
    assert RAM(12487) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12487)))) severity failure;
    assert RAM(12488) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12488)))) severity failure;
    assert RAM(12489) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12489)))) severity failure;
    assert RAM(12490) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12490)))) severity failure;
    assert RAM(12491) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12491)))) severity failure;
    assert RAM(12492) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12492)))) severity failure;
    assert RAM(12493) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12493)))) severity failure;
    assert RAM(12494) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12494)))) severity failure;
    assert RAM(12495) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12495)))) severity failure;
    assert RAM(12496) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12496)))) severity failure;
    assert RAM(12497) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12497)))) severity failure;
    assert RAM(12498) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12498)))) severity failure;
    assert RAM(12499) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12499)))) severity failure;
    assert RAM(12500) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12500)))) severity failure;
    assert RAM(12501) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12501)))) severity failure;
    assert RAM(12502) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12502)))) severity failure;
    assert RAM(12503) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12503)))) severity failure;
    assert RAM(12504) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12504)))) severity failure;
    assert RAM(12505) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12505)))) severity failure;
    assert RAM(12506) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12506)))) severity failure;
    assert RAM(12507) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12507)))) severity failure;
    assert RAM(12508) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12508)))) severity failure;
    assert RAM(12509) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12509)))) severity failure;
    assert RAM(12510) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12510)))) severity failure;
    assert RAM(12511) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12511)))) severity failure;
    assert RAM(12512) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12512)))) severity failure;
    assert RAM(12513) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12513)))) severity failure;
    assert RAM(12514) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12514)))) severity failure;
    assert RAM(12515) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12515)))) severity failure;
    assert RAM(12516) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12516)))) severity failure;
    assert RAM(12517) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12517)))) severity failure;
    assert RAM(12518) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12518)))) severity failure;
    assert RAM(12519) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12519)))) severity failure;
    assert RAM(12520) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12520)))) severity failure;
    assert RAM(12521) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12521)))) severity failure;
    assert RAM(12522) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12522)))) severity failure;
    assert RAM(12523) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12523)))) severity failure;
    assert RAM(12524) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12524)))) severity failure;
    assert RAM(12525) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12525)))) severity failure;
    assert RAM(12526) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12526)))) severity failure;
    assert RAM(12527) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12527)))) severity failure;
    assert RAM(12528) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12528)))) severity failure;
    assert RAM(12529) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12529)))) severity failure;
    assert RAM(12530) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12530)))) severity failure;
    assert RAM(12531) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12531)))) severity failure;
    assert RAM(12532) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12532)))) severity failure;
    assert RAM(12533) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12533)))) severity failure;
    assert RAM(12534) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12534)))) severity failure;
    assert RAM(12535) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12535)))) severity failure;
    assert RAM(12536) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12536)))) severity failure;
    assert RAM(12537) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12537)))) severity failure;
    assert RAM(12538) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12538)))) severity failure;
    assert RAM(12539) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12539)))) severity failure;
    assert RAM(12540) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12540)))) severity failure;
    assert RAM(12541) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12541)))) severity failure;
    assert RAM(12542) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12542)))) severity failure;
    assert RAM(12543) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12543)))) severity failure;
    assert RAM(12544) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12544)))) severity failure;
    assert RAM(12545) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12545)))) severity failure;
    assert RAM(12546) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12546)))) severity failure;
    assert RAM(12547) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12547)))) severity failure;
    assert RAM(12548) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12548)))) severity failure;
    assert RAM(12549) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12549)))) severity failure;
    assert RAM(12550) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12550)))) severity failure;
    assert RAM(12551) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12551)))) severity failure;
    assert RAM(12552) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12552)))) severity failure;
    assert RAM(12553) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12553)))) severity failure;
    assert RAM(12554) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12554)))) severity failure;
    assert RAM(12555) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12555)))) severity failure;
    assert RAM(12556) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12556)))) severity failure;
    assert RAM(12557) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12557)))) severity failure;
    assert RAM(12558) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12558)))) severity failure;
    assert RAM(12559) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12559)))) severity failure;
    assert RAM(12560) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12560)))) severity failure;
    assert RAM(12561) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12561)))) severity failure;
    assert RAM(12562) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12562)))) severity failure;
    assert RAM(12563) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12563)))) severity failure;
    assert RAM(12564) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12564)))) severity failure;
    assert RAM(12565) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12565)))) severity failure;
    assert RAM(12566) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12566)))) severity failure;
    assert RAM(12567) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12567)))) severity failure;
    assert RAM(12568) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12568)))) severity failure;
    assert RAM(12569) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12569)))) severity failure;
    assert RAM(12570) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12570)))) severity failure;
    assert RAM(12571) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12571)))) severity failure;
    assert RAM(12572) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12572)))) severity failure;
    assert RAM(12573) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12573)))) severity failure;
    assert RAM(12574) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12574)))) severity failure;
    assert RAM(12575) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12575)))) severity failure;
    assert RAM(12576) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12576)))) severity failure;
    assert RAM(12577) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12577)))) severity failure;
    assert RAM(12578) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12578)))) severity failure;
    assert RAM(12579) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12579)))) severity failure;
    assert RAM(12580) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12580)))) severity failure;
    assert RAM(12581) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12581)))) severity failure;
    assert RAM(12582) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12582)))) severity failure;
    assert RAM(12583) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12583)))) severity failure;
    assert RAM(12584) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12584)))) severity failure;
    assert RAM(12585) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12585)))) severity failure;
    assert RAM(12586) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12586)))) severity failure;
    assert RAM(12587) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12587)))) severity failure;
    assert RAM(12588) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12588)))) severity failure;
    assert RAM(12589) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12589)))) severity failure;
    assert RAM(12590) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12590)))) severity failure;
    assert RAM(12591) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12591)))) severity failure;
    assert RAM(12592) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12592)))) severity failure;
    assert RAM(12593) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12593)))) severity failure;
    assert RAM(12594) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12594)))) severity failure;
    assert RAM(12595) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12595)))) severity failure;
    assert RAM(12596) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12596)))) severity failure;
    assert RAM(12597) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12597)))) severity failure;
    assert RAM(12598) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12598)))) severity failure;
    assert RAM(12599) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12599)))) severity failure;
    assert RAM(12600) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12600)))) severity failure;
    assert RAM(12601) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12601)))) severity failure;
    assert RAM(12602) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12602)))) severity failure;
    assert RAM(12603) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12603)))) severity failure;
    assert RAM(12604) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12604)))) severity failure;
    assert RAM(12605) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12605)))) severity failure;
    assert RAM(12606) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12606)))) severity failure;
    assert RAM(12607) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12607)))) severity failure;
    assert RAM(12608) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12608)))) severity failure;
    assert RAM(12609) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12609)))) severity failure;
    assert RAM(12610) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12610)))) severity failure;
    assert RAM(12611) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12611)))) severity failure;
    assert RAM(12612) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12612)))) severity failure;
    assert RAM(12613) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12613)))) severity failure;
    assert RAM(12614) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12614)))) severity failure;
    assert RAM(12615) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12615)))) severity failure;
    assert RAM(12616) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12616)))) severity failure;
    assert RAM(12617) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12617)))) severity failure;
    assert RAM(12618) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12618)))) severity failure;
    assert RAM(12619) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12619)))) severity failure;
    assert RAM(12620) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12620)))) severity failure;
    assert RAM(12621) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12621)))) severity failure;
    assert RAM(12622) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12622)))) severity failure;
    assert RAM(12623) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12623)))) severity failure;
    assert RAM(12624) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12624)))) severity failure;
    assert RAM(12625) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12625)))) severity failure;
    assert RAM(12626) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12626)))) severity failure;
    assert RAM(12627) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12627)))) severity failure;
    assert RAM(12628) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12628)))) severity failure;
    assert RAM(12629) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12629)))) severity failure;
    assert RAM(12630) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12630)))) severity failure;
    assert RAM(12631) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12631)))) severity failure;
    assert RAM(12632) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12632)))) severity failure;
    assert RAM(12633) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12633)))) severity failure;
    assert RAM(12634) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12634)))) severity failure;
    assert RAM(12635) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12635)))) severity failure;
    assert RAM(12636) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12636)))) severity failure;
    assert RAM(12637) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12637)))) severity failure;
    assert RAM(12638) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12638)))) severity failure;
    assert RAM(12639) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12639)))) severity failure;
    assert RAM(12640) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12640)))) severity failure;
    assert RAM(12641) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12641)))) severity failure;
    assert RAM(12642) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12642)))) severity failure;
    assert RAM(12643) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12643)))) severity failure;
    assert RAM(12644) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12644)))) severity failure;
    assert RAM(12645) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12645)))) severity failure;
    assert RAM(12646) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12646)))) severity failure;
    assert RAM(12647) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12647)))) severity failure;
    assert RAM(12648) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12648)))) severity failure;
    assert RAM(12649) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12649)))) severity failure;
    assert RAM(12650) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12650)))) severity failure;
    assert RAM(12651) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12651)))) severity failure;
    assert RAM(12652) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12652)))) severity failure;
    assert RAM(12653) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12653)))) severity failure;
    assert RAM(12654) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12654)))) severity failure;
    assert RAM(12655) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12655)))) severity failure;
    assert RAM(12656) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12656)))) severity failure;
    assert RAM(12657) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12657)))) severity failure;
    assert RAM(12658) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12658)))) severity failure;
    assert RAM(12659) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12659)))) severity failure;
    assert RAM(12660) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12660)))) severity failure;
    assert RAM(12661) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12661)))) severity failure;
    assert RAM(12662) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12662)))) severity failure;
    assert RAM(12663) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12663)))) severity failure;
    assert RAM(12664) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12664)))) severity failure;
    assert RAM(12665) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12665)))) severity failure;
    assert RAM(12666) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12666)))) severity failure;
    assert RAM(12667) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12667)))) severity failure;
    assert RAM(12668) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12668)))) severity failure;
    assert RAM(12669) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12669)))) severity failure;
    assert RAM(12670) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12670)))) severity failure;
    assert RAM(12671) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12671)))) severity failure;
    assert RAM(12672) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12672)))) severity failure;
    assert RAM(12673) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12673)))) severity failure;
    assert RAM(12674) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12674)))) severity failure;
    assert RAM(12675) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12675)))) severity failure;
    assert RAM(12676) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12676)))) severity failure;
    assert RAM(12677) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12677)))) severity failure;
    assert RAM(12678) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12678)))) severity failure;
    assert RAM(12679) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12679)))) severity failure;
    assert RAM(12680) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12680)))) severity failure;
    assert RAM(12681) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12681)))) severity failure;
    assert RAM(12682) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12682)))) severity failure;
    assert RAM(12683) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12683)))) severity failure;
    assert RAM(12684) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12684)))) severity failure;
    assert RAM(12685) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12685)))) severity failure;
    assert RAM(12686) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12686)))) severity failure;
    assert RAM(12687) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12687)))) severity failure;
    assert RAM(12688) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12688)))) severity failure;
    assert RAM(12689) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12689)))) severity failure;
    assert RAM(12690) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12690)))) severity failure;
    assert RAM(12691) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12691)))) severity failure;
    assert RAM(12692) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12692)))) severity failure;
    assert RAM(12693) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12693)))) severity failure;
    assert RAM(12694) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12694)))) severity failure;
    assert RAM(12695) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12695)))) severity failure;
    assert RAM(12696) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12696)))) severity failure;
    assert RAM(12697) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12697)))) severity failure;
    assert RAM(12698) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12698)))) severity failure;
    assert RAM(12699) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12699)))) severity failure;
    assert RAM(12700) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12700)))) severity failure;
    assert RAM(12701) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12701)))) severity failure;
    assert RAM(12702) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12702)))) severity failure;
    assert RAM(12703) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12703)))) severity failure;
    assert RAM(12704) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12704)))) severity failure;
    assert RAM(12705) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12705)))) severity failure;
    assert RAM(12706) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12706)))) severity failure;
    assert RAM(12707) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12707)))) severity failure;
    assert RAM(12708) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12708)))) severity failure;
    assert RAM(12709) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12709)))) severity failure;
    assert RAM(12710) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12710)))) severity failure;
    assert RAM(12711) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12711)))) severity failure;
    assert RAM(12712) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12712)))) severity failure;
    assert RAM(12713) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12713)))) severity failure;
    assert RAM(12714) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12714)))) severity failure;
    assert RAM(12715) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12715)))) severity failure;
    assert RAM(12716) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12716)))) severity failure;
    assert RAM(12717) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12717)))) severity failure;
    assert RAM(12718) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12718)))) severity failure;
    assert RAM(12719) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12719)))) severity failure;
    assert RAM(12720) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12720)))) severity failure;
    assert RAM(12721) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12721)))) severity failure;
    assert RAM(12722) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12722)))) severity failure;
    assert RAM(12723) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12723)))) severity failure;
    assert RAM(12724) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12724)))) severity failure;
    assert RAM(12725) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12725)))) severity failure;
    assert RAM(12726) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12726)))) severity failure;
    assert RAM(12727) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12727)))) severity failure;
    assert RAM(12728) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12728)))) severity failure;
    assert RAM(12729) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12729)))) severity failure;
    assert RAM(12730) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12730)))) severity failure;
    assert RAM(12731) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12731)))) severity failure;
    assert RAM(12732) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12732)))) severity failure;
    assert RAM(12733) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12733)))) severity failure;
    assert RAM(12734) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12734)))) severity failure;
    assert RAM(12735) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12735)))) severity failure;
    assert RAM(12736) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12736)))) severity failure;
    assert RAM(12737) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12737)))) severity failure;
    assert RAM(12738) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12738)))) severity failure;
    assert RAM(12739) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12739)))) severity failure;
    assert RAM(12740) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12740)))) severity failure;
    assert RAM(12741) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12741)))) severity failure;
    assert RAM(12742) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12742)))) severity failure;
    assert RAM(12743) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12743)))) severity failure;
    assert RAM(12744) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12744)))) severity failure;
    assert RAM(12745) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12745)))) severity failure;
    assert RAM(12746) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12746)))) severity failure;
    assert RAM(12747) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12747)))) severity failure;
    assert RAM(12748) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12748)))) severity failure;
    assert RAM(12749) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12749)))) severity failure;
    assert RAM(12750) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12750)))) severity failure;
    assert RAM(12751) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12751)))) severity failure;
    assert RAM(12752) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12752)))) severity failure;
    assert RAM(12753) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12753)))) severity failure;
    assert RAM(12754) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12754)))) severity failure;
    assert RAM(12755) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12755)))) severity failure;
    assert RAM(12756) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12756)))) severity failure;
    assert RAM(12757) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12757)))) severity failure;
    assert RAM(12758) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12758)))) severity failure;
    assert RAM(12759) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12759)))) severity failure;
    assert RAM(12760) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12760)))) severity failure;
    assert RAM(12761) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12761)))) severity failure;
    assert RAM(12762) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12762)))) severity failure;
    assert RAM(12763) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12763)))) severity failure;
    assert RAM(12764) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12764)))) severity failure;
    assert RAM(12765) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12765)))) severity failure;
    assert RAM(12766) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12766)))) severity failure;
    assert RAM(12767) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12767)))) severity failure;
    assert RAM(12768) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12768)))) severity failure;
    assert RAM(12769) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12769)))) severity failure;
    assert RAM(12770) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12770)))) severity failure;
    assert RAM(12771) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12771)))) severity failure;
    assert RAM(12772) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12772)))) severity failure;
    assert RAM(12773) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12773)))) severity failure;
    assert RAM(12774) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12774)))) severity failure;
    assert RAM(12775) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12775)))) severity failure;
    assert RAM(12776) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12776)))) severity failure;
    assert RAM(12777) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12777)))) severity failure;
    assert RAM(12778) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12778)))) severity failure;
    assert RAM(12779) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12779)))) severity failure;
    assert RAM(12780) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12780)))) severity failure;
    assert RAM(12781) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12781)))) severity failure;
    assert RAM(12782) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12782)))) severity failure;
    assert RAM(12783) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12783)))) severity failure;
    assert RAM(12784) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12784)))) severity failure;
    assert RAM(12785) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12785)))) severity failure;
    assert RAM(12786) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12786)))) severity failure;
    assert RAM(12787) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12787)))) severity failure;
    assert RAM(12788) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12788)))) severity failure;
    assert RAM(12789) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12789)))) severity failure;
    assert RAM(12790) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12790)))) severity failure;
    assert RAM(12791) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12791)))) severity failure;
    assert RAM(12792) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12792)))) severity failure;
    assert RAM(12793) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12793)))) severity failure;
    assert RAM(12794) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12794)))) severity failure;
    assert RAM(12795) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12795)))) severity failure;
    assert RAM(12796) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12796)))) severity failure;
    assert RAM(12797) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12797)))) severity failure;
    assert RAM(12798) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12798)))) severity failure;
    assert RAM(12799) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12799)))) severity failure;
    assert RAM(12800) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12800)))) severity failure;
    assert RAM(12801) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12801)))) severity failure;
    assert RAM(12802) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12802)))) severity failure;
    assert RAM(12803) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12803)))) severity failure;
    assert RAM(12804) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12804)))) severity failure;
    assert RAM(12805) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12805)))) severity failure;
    assert RAM(12806) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12806)))) severity failure;
    assert RAM(12807) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12807)))) severity failure;
    assert RAM(12808) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12808)))) severity failure;
    assert RAM(12809) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12809)))) severity failure;
    assert RAM(12810) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12810)))) severity failure;
    assert RAM(12811) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12811)))) severity failure;
    assert RAM(12812) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12812)))) severity failure;
    assert RAM(12813) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12813)))) severity failure;
    assert RAM(12814) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12814)))) severity failure;
    assert RAM(12815) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12815)))) severity failure;
    assert RAM(12816) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12816)))) severity failure;
    assert RAM(12817) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12817)))) severity failure;
    assert RAM(12818) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12818)))) severity failure;
    assert RAM(12819) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12819)))) severity failure;
    assert RAM(12820) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12820)))) severity failure;
    assert RAM(12821) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12821)))) severity failure;
    assert RAM(12822) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12822)))) severity failure;
    assert RAM(12823) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12823)))) severity failure;
    assert RAM(12824) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12824)))) severity failure;
    assert RAM(12825) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12825)))) severity failure;
    assert RAM(12826) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12826)))) severity failure;
    assert RAM(12827) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12827)))) severity failure;
    assert RAM(12828) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12828)))) severity failure;
    assert RAM(12829) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12829)))) severity failure;
    assert RAM(12830) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12830)))) severity failure;
    assert RAM(12831) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12831)))) severity failure;
    assert RAM(12832) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12832)))) severity failure;
    assert RAM(12833) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12833)))) severity failure;
    assert RAM(12834) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12834)))) severity failure;
    assert RAM(12835) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12835)))) severity failure;
    assert RAM(12836) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12836)))) severity failure;
    assert RAM(12837) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12837)))) severity failure;
    assert RAM(12838) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12838)))) severity failure;
    assert RAM(12839) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12839)))) severity failure;
    assert RAM(12840) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12840)))) severity failure;
    assert RAM(12841) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12841)))) severity failure;
    assert RAM(12842) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12842)))) severity failure;
    assert RAM(12843) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12843)))) severity failure;
    assert RAM(12844) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12844)))) severity failure;
    assert RAM(12845) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12845)))) severity failure;
    assert RAM(12846) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12846)))) severity failure;
    assert RAM(12847) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12847)))) severity failure;
    assert RAM(12848) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12848)))) severity failure;
    assert RAM(12849) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12849)))) severity failure;
    assert RAM(12850) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12850)))) severity failure;
    assert RAM(12851) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12851)))) severity failure;
    assert RAM(12852) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12852)))) severity failure;
    assert RAM(12853) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12853)))) severity failure;
    assert RAM(12854) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12854)))) severity failure;
    assert RAM(12855) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12855)))) severity failure;
    assert RAM(12856) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12856)))) severity failure;
    assert RAM(12857) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12857)))) severity failure;
    assert RAM(12858) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12858)))) severity failure;
    assert RAM(12859) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12859)))) severity failure;
    assert RAM(12860) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12860)))) severity failure;
    assert RAM(12861) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12861)))) severity failure;
    assert RAM(12862) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12862)))) severity failure;
    assert RAM(12863) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12863)))) severity failure;
    assert RAM(12864) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12864)))) severity failure;
    assert RAM(12865) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12865)))) severity failure;
    assert RAM(12866) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12866)))) severity failure;
    assert RAM(12867) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12867)))) severity failure;
    assert RAM(12868) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12868)))) severity failure;
    assert RAM(12869) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12869)))) severity failure;
    assert RAM(12870) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12870)))) severity failure;
    assert RAM(12871) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12871)))) severity failure;
    assert RAM(12872) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12872)))) severity failure;
    assert RAM(12873) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12873)))) severity failure;
    assert RAM(12874) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12874)))) severity failure;
    assert RAM(12875) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12875)))) severity failure;
    assert RAM(12876) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12876)))) severity failure;
    assert RAM(12877) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12877)))) severity failure;
    assert RAM(12878) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12878)))) severity failure;
    assert RAM(12879) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12879)))) severity failure;
    assert RAM(12880) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12880)))) severity failure;
    assert RAM(12881) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12881)))) severity failure;
    assert RAM(12882) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12882)))) severity failure;
    assert RAM(12883) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12883)))) severity failure;
    assert RAM(12884) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12884)))) severity failure;
    assert RAM(12885) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12885)))) severity failure;
    assert RAM(12886) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12886)))) severity failure;
    assert RAM(12887) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12887)))) severity failure;
    assert RAM(12888) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12888)))) severity failure;
    assert RAM(12889) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12889)))) severity failure;
    assert RAM(12890) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12890)))) severity failure;
    assert RAM(12891) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12891)))) severity failure;
    assert RAM(12892) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12892)))) severity failure;
    assert RAM(12893) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12893)))) severity failure;
    assert RAM(12894) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12894)))) severity failure;
    assert RAM(12895) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12895)))) severity failure;
    assert RAM(12896) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12896)))) severity failure;
    assert RAM(12897) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12897)))) severity failure;
    assert RAM(12898) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12898)))) severity failure;
    assert RAM(12899) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12899)))) severity failure;
    assert RAM(12900) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12900)))) severity failure;
    assert RAM(12901) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12901)))) severity failure;
    assert RAM(12902) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12902)))) severity failure;
    assert RAM(12903) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12903)))) severity failure;
    assert RAM(12904) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12904)))) severity failure;
    assert RAM(12905) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12905)))) severity failure;
    assert RAM(12906) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12906)))) severity failure;
    assert RAM(12907) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12907)))) severity failure;
    assert RAM(12908) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12908)))) severity failure;
    assert RAM(12909) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12909)))) severity failure;
    assert RAM(12910) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12910)))) severity failure;
    assert RAM(12911) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12911)))) severity failure;
    assert RAM(12912) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12912)))) severity failure;
    assert RAM(12913) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12913)))) severity failure;
    assert RAM(12914) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12914)))) severity failure;
    assert RAM(12915) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12915)))) severity failure;
    assert RAM(12916) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12916)))) severity failure;
    assert RAM(12917) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12917)))) severity failure;
    assert RAM(12918) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12918)))) severity failure;
    assert RAM(12919) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12919)))) severity failure;
    assert RAM(12920) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12920)))) severity failure;
    assert RAM(12921) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12921)))) severity failure;
    assert RAM(12922) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12922)))) severity failure;
    assert RAM(12923) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12923)))) severity failure;
    assert RAM(12924) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12924)))) severity failure;
    assert RAM(12925) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12925)))) severity failure;
    assert RAM(12926) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12926)))) severity failure;
    assert RAM(12927) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12927)))) severity failure;
    assert RAM(12928) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12928)))) severity failure;
    assert RAM(12929) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12929)))) severity failure;
    assert RAM(12930) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12930)))) severity failure;
    assert RAM(12931) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12931)))) severity failure;
    assert RAM(12932) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12932)))) severity failure;
    assert RAM(12933) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12933)))) severity failure;
    assert RAM(12934) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12934)))) severity failure;
    assert RAM(12935) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12935)))) severity failure;
    assert RAM(12936) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12936)))) severity failure;
    assert RAM(12937) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12937)))) severity failure;
    assert RAM(12938) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12938)))) severity failure;
    assert RAM(12939) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12939)))) severity failure;
    assert RAM(12940) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12940)))) severity failure;
    assert RAM(12941) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12941)))) severity failure;
    assert RAM(12942) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12942)))) severity failure;
    assert RAM(12943) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12943)))) severity failure;
    assert RAM(12944) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12944)))) severity failure;
    assert RAM(12945) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12945)))) severity failure;
    assert RAM(12946) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12946)))) severity failure;
    assert RAM(12947) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12947)))) severity failure;
    assert RAM(12948) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12948)))) severity failure;
    assert RAM(12949) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12949)))) severity failure;
    assert RAM(12950) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12950)))) severity failure;
    assert RAM(12951) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12951)))) severity failure;
    assert RAM(12952) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12952)))) severity failure;
    assert RAM(12953) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12953)))) severity failure;
    assert RAM(12954) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12954)))) severity failure;
    assert RAM(12955) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12955)))) severity failure;
    assert RAM(12956) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12956)))) severity failure;
    assert RAM(12957) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12957)))) severity failure;
    assert RAM(12958) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12958)))) severity failure;
    assert RAM(12959) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12959)))) severity failure;
    assert RAM(12960) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12960)))) severity failure;
    assert RAM(12961) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12961)))) severity failure;
    assert RAM(12962) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12962)))) severity failure;
    assert RAM(12963) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12963)))) severity failure;
    assert RAM(12964) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12964)))) severity failure;
    assert RAM(12965) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12965)))) severity failure;
    assert RAM(12966) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12966)))) severity failure;
    assert RAM(12967) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12967)))) severity failure;
    assert RAM(12968) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12968)))) severity failure;
    assert RAM(12969) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12969)))) severity failure;
    assert RAM(12970) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12970)))) severity failure;
    assert RAM(12971) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12971)))) severity failure;
    assert RAM(12972) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12972)))) severity failure;
    assert RAM(12973) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12973)))) severity failure;
    assert RAM(12974) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12974)))) severity failure;
    assert RAM(12975) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12975)))) severity failure;
    assert RAM(12976) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12976)))) severity failure;
    assert RAM(12977) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12977)))) severity failure;
    assert RAM(12978) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12978)))) severity failure;
    assert RAM(12979) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12979)))) severity failure;
    assert RAM(12980) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12980)))) severity failure;
    assert RAM(12981) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12981)))) severity failure;
    assert RAM(12982) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12982)))) severity failure;
    assert RAM(12983) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12983)))) severity failure;
    assert RAM(12984) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12984)))) severity failure;
    assert RAM(12985) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12985)))) severity failure;
    assert RAM(12986) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12986)))) severity failure;
    assert RAM(12987) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12987)))) severity failure;
    assert RAM(12988) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12988)))) severity failure;
    assert RAM(12989) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12989)))) severity failure;
    assert RAM(12990) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12990)))) severity failure;
    assert RAM(12991) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12991)))) severity failure;
    assert RAM(12992) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12992)))) severity failure;
    assert RAM(12993) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12993)))) severity failure;
    assert RAM(12994) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12994)))) severity failure;
    assert RAM(12995) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12995)))) severity failure;
    assert RAM(12996) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(12996)))) severity failure;
    assert RAM(12997) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12997)))) severity failure;
    assert RAM(12998) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12998)))) severity failure;
    assert RAM(12999) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(12999)))) severity failure;
    assert RAM(13000) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13000)))) severity failure;
    assert RAM(13001) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13001)))) severity failure;
    assert RAM(13002) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13002)))) severity failure;
    assert RAM(13003) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13003)))) severity failure;
    assert RAM(13004) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13004)))) severity failure;
    assert RAM(13005) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13005)))) severity failure;
    assert RAM(13006) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13006)))) severity failure;
    assert RAM(13007) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13007)))) severity failure;
    assert RAM(13008) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13008)))) severity failure;
    assert RAM(13009) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13009)))) severity failure;
    assert RAM(13010) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13010)))) severity failure;
    assert RAM(13011) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13011)))) severity failure;
    assert RAM(13012) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13012)))) severity failure;
    assert RAM(13013) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13013)))) severity failure;
    assert RAM(13014) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13014)))) severity failure;
    assert RAM(13015) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13015)))) severity failure;
    assert RAM(13016) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13016)))) severity failure;
    assert RAM(13017) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13017)))) severity failure;
    assert RAM(13018) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13018)))) severity failure;
    assert RAM(13019) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13019)))) severity failure;
    assert RAM(13020) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13020)))) severity failure;
    assert RAM(13021) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13021)))) severity failure;
    assert RAM(13022) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13022)))) severity failure;
    assert RAM(13023) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13023)))) severity failure;
    assert RAM(13024) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13024)))) severity failure;
    assert RAM(13025) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13025)))) severity failure;
    assert RAM(13026) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13026)))) severity failure;
    assert RAM(13027) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13027)))) severity failure;
    assert RAM(13028) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13028)))) severity failure;
    assert RAM(13029) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13029)))) severity failure;
    assert RAM(13030) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13030)))) severity failure;
    assert RAM(13031) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13031)))) severity failure;
    assert RAM(13032) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13032)))) severity failure;
    assert RAM(13033) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13033)))) severity failure;
    assert RAM(13034) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13034)))) severity failure;
    assert RAM(13035) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13035)))) severity failure;
    assert RAM(13036) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13036)))) severity failure;
    assert RAM(13037) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13037)))) severity failure;
    assert RAM(13038) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13038)))) severity failure;
    assert RAM(13039) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13039)))) severity failure;
    assert RAM(13040) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13040)))) severity failure;
    assert RAM(13041) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13041)))) severity failure;
    assert RAM(13042) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13042)))) severity failure;
    assert RAM(13043) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13043)))) severity failure;
    assert RAM(13044) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13044)))) severity failure;
    assert RAM(13045) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13045)))) severity failure;
    assert RAM(13046) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13046)))) severity failure;
    assert RAM(13047) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13047)))) severity failure;
    assert RAM(13048) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13048)))) severity failure;
    assert RAM(13049) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13049)))) severity failure;
    assert RAM(13050) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13050)))) severity failure;
    assert RAM(13051) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13051)))) severity failure;
    assert RAM(13052) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13052)))) severity failure;
    assert RAM(13053) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13053)))) severity failure;
    assert RAM(13054) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13054)))) severity failure;
    assert RAM(13055) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13055)))) severity failure;
    assert RAM(13056) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13056)))) severity failure;
    assert RAM(13057) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13057)))) severity failure;
    assert RAM(13058) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13058)))) severity failure;
    assert RAM(13059) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13059)))) severity failure;
    assert RAM(13060) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13060)))) severity failure;
    assert RAM(13061) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13061)))) severity failure;
    assert RAM(13062) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13062)))) severity failure;
    assert RAM(13063) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13063)))) severity failure;
    assert RAM(13064) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13064)))) severity failure;
    assert RAM(13065) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13065)))) severity failure;
    assert RAM(13066) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13066)))) severity failure;
    assert RAM(13067) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13067)))) severity failure;
    assert RAM(13068) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13068)))) severity failure;
    assert RAM(13069) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13069)))) severity failure;
    assert RAM(13070) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13070)))) severity failure;
    assert RAM(13071) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13071)))) severity failure;
    assert RAM(13072) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13072)))) severity failure;
    assert RAM(13073) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13073)))) severity failure;
    assert RAM(13074) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13074)))) severity failure;
    assert RAM(13075) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13075)))) severity failure;
    assert RAM(13076) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13076)))) severity failure;
    assert RAM(13077) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13077)))) severity failure;
    assert RAM(13078) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13078)))) severity failure;
    assert RAM(13079) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13079)))) severity failure;
    assert RAM(13080) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13080)))) severity failure;
    assert RAM(13081) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13081)))) severity failure;
    assert RAM(13082) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13082)))) severity failure;
    assert RAM(13083) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13083)))) severity failure;
    assert RAM(13084) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13084)))) severity failure;
    assert RAM(13085) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13085)))) severity failure;
    assert RAM(13086) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13086)))) severity failure;
    assert RAM(13087) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13087)))) severity failure;
    assert RAM(13088) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13088)))) severity failure;
    assert RAM(13089) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13089)))) severity failure;
    assert RAM(13090) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13090)))) severity failure;
    assert RAM(13091) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13091)))) severity failure;
    assert RAM(13092) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13092)))) severity failure;
    assert RAM(13093) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13093)))) severity failure;
    assert RAM(13094) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13094)))) severity failure;
    assert RAM(13095) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13095)))) severity failure;
    assert RAM(13096) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13096)))) severity failure;
    assert RAM(13097) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13097)))) severity failure;
    assert RAM(13098) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13098)))) severity failure;
    assert RAM(13099) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13099)))) severity failure;
    assert RAM(13100) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13100)))) severity failure;
    assert RAM(13101) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13101)))) severity failure;
    assert RAM(13102) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13102)))) severity failure;
    assert RAM(13103) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13103)))) severity failure;
    assert RAM(13104) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13104)))) severity failure;
    assert RAM(13105) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13105)))) severity failure;
    assert RAM(13106) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13106)))) severity failure;
    assert RAM(13107) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13107)))) severity failure;
    assert RAM(13108) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13108)))) severity failure;
    assert RAM(13109) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13109)))) severity failure;
    assert RAM(13110) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13110)))) severity failure;
    assert RAM(13111) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13111)))) severity failure;
    assert RAM(13112) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13112)))) severity failure;
    assert RAM(13113) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13113)))) severity failure;
    assert RAM(13114) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13114)))) severity failure;
    assert RAM(13115) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13115)))) severity failure;
    assert RAM(13116) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13116)))) severity failure;
    assert RAM(13117) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13117)))) severity failure;
    assert RAM(13118) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13118)))) severity failure;
    assert RAM(13119) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13119)))) severity failure;
    assert RAM(13120) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13120)))) severity failure;
    assert RAM(13121) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13121)))) severity failure;
    assert RAM(13122) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13122)))) severity failure;
    assert RAM(13123) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13123)))) severity failure;
    assert RAM(13124) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13124)))) severity failure;
    assert RAM(13125) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13125)))) severity failure;
    assert RAM(13126) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13126)))) severity failure;
    assert RAM(13127) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13127)))) severity failure;
    assert RAM(13128) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13128)))) severity failure;
    assert RAM(13129) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13129)))) severity failure;
    assert RAM(13130) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13130)))) severity failure;
    assert RAM(13131) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13131)))) severity failure;
    assert RAM(13132) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13132)))) severity failure;
    assert RAM(13133) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13133)))) severity failure;
    assert RAM(13134) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13134)))) severity failure;
    assert RAM(13135) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13135)))) severity failure;
    assert RAM(13136) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13136)))) severity failure;
    assert RAM(13137) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13137)))) severity failure;
    assert RAM(13138) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13138)))) severity failure;
    assert RAM(13139) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13139)))) severity failure;
    assert RAM(13140) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13140)))) severity failure;
    assert RAM(13141) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13141)))) severity failure;
    assert RAM(13142) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13142)))) severity failure;
    assert RAM(13143) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13143)))) severity failure;
    assert RAM(13144) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13144)))) severity failure;
    assert RAM(13145) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13145)))) severity failure;
    assert RAM(13146) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13146)))) severity failure;
    assert RAM(13147) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13147)))) severity failure;
    assert RAM(13148) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13148)))) severity failure;
    assert RAM(13149) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13149)))) severity failure;
    assert RAM(13150) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13150)))) severity failure;
    assert RAM(13151) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13151)))) severity failure;
    assert RAM(13152) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13152)))) severity failure;
    assert RAM(13153) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13153)))) severity failure;
    assert RAM(13154) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13154)))) severity failure;
    assert RAM(13155) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13155)))) severity failure;
    assert RAM(13156) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13156)))) severity failure;
    assert RAM(13157) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13157)))) severity failure;
    assert RAM(13158) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13158)))) severity failure;
    assert RAM(13159) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13159)))) severity failure;
    assert RAM(13160) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13160)))) severity failure;
    assert RAM(13161) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13161)))) severity failure;
    assert RAM(13162) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13162)))) severity failure;
    assert RAM(13163) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13163)))) severity failure;
    assert RAM(13164) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13164)))) severity failure;
    assert RAM(13165) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13165)))) severity failure;
    assert RAM(13166) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13166)))) severity failure;
    assert RAM(13167) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13167)))) severity failure;
    assert RAM(13168) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13168)))) severity failure;
    assert RAM(13169) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13169)))) severity failure;
    assert RAM(13170) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13170)))) severity failure;
    assert RAM(13171) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13171)))) severity failure;
    assert RAM(13172) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13172)))) severity failure;
    assert RAM(13173) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13173)))) severity failure;
    assert RAM(13174) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13174)))) severity failure;
    assert RAM(13175) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13175)))) severity failure;
    assert RAM(13176) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13176)))) severity failure;
    assert RAM(13177) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13177)))) severity failure;
    assert RAM(13178) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13178)))) severity failure;
    assert RAM(13179) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13179)))) severity failure;
    assert RAM(13180) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13180)))) severity failure;
    assert RAM(13181) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13181)))) severity failure;
    assert RAM(13182) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13182)))) severity failure;
    assert RAM(13183) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13183)))) severity failure;
    assert RAM(13184) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13184)))) severity failure;
    assert RAM(13185) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13185)))) severity failure;
    assert RAM(13186) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13186)))) severity failure;
    assert RAM(13187) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13187)))) severity failure;
    assert RAM(13188) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13188)))) severity failure;
    assert RAM(13189) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13189)))) severity failure;
    assert RAM(13190) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13190)))) severity failure;
    assert RAM(13191) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13191)))) severity failure;
    assert RAM(13192) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13192)))) severity failure;
    assert RAM(13193) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13193)))) severity failure;
    assert RAM(13194) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13194)))) severity failure;
    assert RAM(13195) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13195)))) severity failure;
    assert RAM(13196) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13196)))) severity failure;
    assert RAM(13197) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13197)))) severity failure;
    assert RAM(13198) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13198)))) severity failure;
    assert RAM(13199) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13199)))) severity failure;
    assert RAM(13200) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13200)))) severity failure;
    assert RAM(13201) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13201)))) severity failure;
    assert RAM(13202) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13202)))) severity failure;
    assert RAM(13203) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13203)))) severity failure;
    assert RAM(13204) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13204)))) severity failure;
    assert RAM(13205) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13205)))) severity failure;
    assert RAM(13206) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13206)))) severity failure;
    assert RAM(13207) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13207)))) severity failure;
    assert RAM(13208) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13208)))) severity failure;
    assert RAM(13209) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13209)))) severity failure;
    assert RAM(13210) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13210)))) severity failure;
    assert RAM(13211) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13211)))) severity failure;
    assert RAM(13212) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13212)))) severity failure;
    assert RAM(13213) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13213)))) severity failure;
    assert RAM(13214) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13214)))) severity failure;
    assert RAM(13215) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13215)))) severity failure;
    assert RAM(13216) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13216)))) severity failure;
    assert RAM(13217) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13217)))) severity failure;
    assert RAM(13218) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13218)))) severity failure;
    assert RAM(13219) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13219)))) severity failure;
    assert RAM(13220) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13220)))) severity failure;
    assert RAM(13221) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13221)))) severity failure;
    assert RAM(13222) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13222)))) severity failure;
    assert RAM(13223) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13223)))) severity failure;
    assert RAM(13224) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13224)))) severity failure;
    assert RAM(13225) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13225)))) severity failure;
    assert RAM(13226) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13226)))) severity failure;
    assert RAM(13227) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13227)))) severity failure;
    assert RAM(13228) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13228)))) severity failure;
    assert RAM(13229) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13229)))) severity failure;
    assert RAM(13230) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13230)))) severity failure;
    assert RAM(13231) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13231)))) severity failure;
    assert RAM(13232) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13232)))) severity failure;
    assert RAM(13233) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13233)))) severity failure;
    assert RAM(13234) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13234)))) severity failure;
    assert RAM(13235) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13235)))) severity failure;
    assert RAM(13236) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13236)))) severity failure;
    assert RAM(13237) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13237)))) severity failure;
    assert RAM(13238) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13238)))) severity failure;
    assert RAM(13239) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13239)))) severity failure;
    assert RAM(13240) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13240)))) severity failure;
    assert RAM(13241) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13241)))) severity failure;
    assert RAM(13242) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13242)))) severity failure;
    assert RAM(13243) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13243)))) severity failure;
    assert RAM(13244) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13244)))) severity failure;
    assert RAM(13245) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13245)))) severity failure;
    assert RAM(13246) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13246)))) severity failure;
    assert RAM(13247) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13247)))) severity failure;
    assert RAM(13248) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13248)))) severity failure;
    assert RAM(13249) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13249)))) severity failure;
    assert RAM(13250) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13250)))) severity failure;
    assert RAM(13251) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13251)))) severity failure;
    assert RAM(13252) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13252)))) severity failure;
    assert RAM(13253) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13253)))) severity failure;
    assert RAM(13254) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13254)))) severity failure;
    assert RAM(13255) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13255)))) severity failure;
    assert RAM(13256) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13256)))) severity failure;
    assert RAM(13257) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13257)))) severity failure;
    assert RAM(13258) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13258)))) severity failure;
    assert RAM(13259) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13259)))) severity failure;
    assert RAM(13260) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13260)))) severity failure;
    assert RAM(13261) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13261)))) severity failure;
    assert RAM(13262) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13262)))) severity failure;
    assert RAM(13263) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13263)))) severity failure;
    assert RAM(13264) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13264)))) severity failure;
    assert RAM(13265) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13265)))) severity failure;
    assert RAM(13266) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13266)))) severity failure;
    assert RAM(13267) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13267)))) severity failure;
    assert RAM(13268) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13268)))) severity failure;
    assert RAM(13269) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13269)))) severity failure;
    assert RAM(13270) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13270)))) severity failure;
    assert RAM(13271) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13271)))) severity failure;
    assert RAM(13272) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13272)))) severity failure;
    assert RAM(13273) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13273)))) severity failure;
    assert RAM(13274) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13274)))) severity failure;
    assert RAM(13275) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13275)))) severity failure;
    assert RAM(13276) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13276)))) severity failure;
    assert RAM(13277) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13277)))) severity failure;
    assert RAM(13278) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13278)))) severity failure;
    assert RAM(13279) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13279)))) severity failure;
    assert RAM(13280) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13280)))) severity failure;
    assert RAM(13281) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13281)))) severity failure;
    assert RAM(13282) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13282)))) severity failure;
    assert RAM(13283) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13283)))) severity failure;
    assert RAM(13284) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13284)))) severity failure;
    assert RAM(13285) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13285)))) severity failure;
    assert RAM(13286) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13286)))) severity failure;
    assert RAM(13287) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13287)))) severity failure;
    assert RAM(13288) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13288)))) severity failure;
    assert RAM(13289) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13289)))) severity failure;
    assert RAM(13290) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13290)))) severity failure;
    assert RAM(13291) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13291)))) severity failure;
    assert RAM(13292) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13292)))) severity failure;
    assert RAM(13293) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13293)))) severity failure;
    assert RAM(13294) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13294)))) severity failure;
    assert RAM(13295) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13295)))) severity failure;
    assert RAM(13296) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13296)))) severity failure;
    assert RAM(13297) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13297)))) severity failure;
    assert RAM(13298) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13298)))) severity failure;
    assert RAM(13299) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13299)))) severity failure;
    assert RAM(13300) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13300)))) severity failure;
    assert RAM(13301) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13301)))) severity failure;
    assert RAM(13302) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13302)))) severity failure;
    assert RAM(13303) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13303)))) severity failure;
    assert RAM(13304) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13304)))) severity failure;
    assert RAM(13305) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13305)))) severity failure;
    assert RAM(13306) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13306)))) severity failure;
    assert RAM(13307) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13307)))) severity failure;
    assert RAM(13308) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13308)))) severity failure;
    assert RAM(13309) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13309)))) severity failure;
    assert RAM(13310) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13310)))) severity failure;
    assert RAM(13311) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13311)))) severity failure;
    assert RAM(13312) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13312)))) severity failure;
    assert RAM(13313) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13313)))) severity failure;
    assert RAM(13314) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13314)))) severity failure;
    assert RAM(13315) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13315)))) severity failure;
    assert RAM(13316) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13316)))) severity failure;
    assert RAM(13317) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13317)))) severity failure;
    assert RAM(13318) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13318)))) severity failure;
    assert RAM(13319) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13319)))) severity failure;
    assert RAM(13320) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13320)))) severity failure;
    assert RAM(13321) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13321)))) severity failure;
    assert RAM(13322) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13322)))) severity failure;
    assert RAM(13323) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13323)))) severity failure;
    assert RAM(13324) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13324)))) severity failure;
    assert RAM(13325) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13325)))) severity failure;
    assert RAM(13326) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13326)))) severity failure;
    assert RAM(13327) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13327)))) severity failure;
    assert RAM(13328) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13328)))) severity failure;
    assert RAM(13329) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13329)))) severity failure;
    assert RAM(13330) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13330)))) severity failure;
    assert RAM(13331) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13331)))) severity failure;
    assert RAM(13332) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13332)))) severity failure;
    assert RAM(13333) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13333)))) severity failure;
    assert RAM(13334) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13334)))) severity failure;
    assert RAM(13335) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13335)))) severity failure;
    assert RAM(13336) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13336)))) severity failure;
    assert RAM(13337) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13337)))) severity failure;
    assert RAM(13338) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13338)))) severity failure;
    assert RAM(13339) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13339)))) severity failure;
    assert RAM(13340) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13340)))) severity failure;
    assert RAM(13341) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13341)))) severity failure;
    assert RAM(13342) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13342)))) severity failure;
    assert RAM(13343) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13343)))) severity failure;
    assert RAM(13344) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13344)))) severity failure;
    assert RAM(13345) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13345)))) severity failure;
    assert RAM(13346) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13346)))) severity failure;
    assert RAM(13347) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13347)))) severity failure;
    assert RAM(13348) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13348)))) severity failure;
    assert RAM(13349) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13349)))) severity failure;
    assert RAM(13350) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13350)))) severity failure;
    assert RAM(13351) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13351)))) severity failure;
    assert RAM(13352) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13352)))) severity failure;
    assert RAM(13353) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13353)))) severity failure;
    assert RAM(13354) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13354)))) severity failure;
    assert RAM(13355) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13355)))) severity failure;
    assert RAM(13356) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13356)))) severity failure;
    assert RAM(13357) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13357)))) severity failure;
    assert RAM(13358) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13358)))) severity failure;
    assert RAM(13359) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13359)))) severity failure;
    assert RAM(13360) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13360)))) severity failure;
    assert RAM(13361) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13361)))) severity failure;
    assert RAM(13362) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13362)))) severity failure;
    assert RAM(13363) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13363)))) severity failure;
    assert RAM(13364) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13364)))) severity failure;
    assert RAM(13365) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13365)))) severity failure;
    assert RAM(13366) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13366)))) severity failure;
    assert RAM(13367) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13367)))) severity failure;
    assert RAM(13368) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13368)))) severity failure;
    assert RAM(13369) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13369)))) severity failure;
    assert RAM(13370) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13370)))) severity failure;
    assert RAM(13371) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13371)))) severity failure;
    assert RAM(13372) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13372)))) severity failure;
    assert RAM(13373) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13373)))) severity failure;
    assert RAM(13374) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13374)))) severity failure;
    assert RAM(13375) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13375)))) severity failure;
    assert RAM(13376) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13376)))) severity failure;
    assert RAM(13377) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13377)))) severity failure;
    assert RAM(13378) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13378)))) severity failure;
    assert RAM(13379) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13379)))) severity failure;
    assert RAM(13380) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13380)))) severity failure;
    assert RAM(13381) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13381)))) severity failure;
    assert RAM(13382) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13382)))) severity failure;
    assert RAM(13383) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13383)))) severity failure;
    assert RAM(13384) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13384)))) severity failure;
    assert RAM(13385) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13385)))) severity failure;
    assert RAM(13386) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13386)))) severity failure;
    assert RAM(13387) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13387)))) severity failure;
    assert RAM(13388) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13388)))) severity failure;
    assert RAM(13389) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13389)))) severity failure;
    assert RAM(13390) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13390)))) severity failure;
    assert RAM(13391) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13391)))) severity failure;
    assert RAM(13392) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13392)))) severity failure;
    assert RAM(13393) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13393)))) severity failure;
    assert RAM(13394) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13394)))) severity failure;
    assert RAM(13395) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13395)))) severity failure;
    assert RAM(13396) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13396)))) severity failure;
    assert RAM(13397) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13397)))) severity failure;
    assert RAM(13398) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13398)))) severity failure;
    assert RAM(13399) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13399)))) severity failure;
    assert RAM(13400) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13400)))) severity failure;
    assert RAM(13401) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13401)))) severity failure;
    assert RAM(13402) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13402)))) severity failure;
    assert RAM(13403) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13403)))) severity failure;
    assert RAM(13404) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13404)))) severity failure;
    assert RAM(13405) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13405)))) severity failure;
    assert RAM(13406) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13406)))) severity failure;
    assert RAM(13407) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13407)))) severity failure;
    assert RAM(13408) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13408)))) severity failure;
    assert RAM(13409) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13409)))) severity failure;
    assert RAM(13410) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13410)))) severity failure;
    assert RAM(13411) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13411)))) severity failure;
    assert RAM(13412) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13412)))) severity failure;
    assert RAM(13413) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13413)))) severity failure;
    assert RAM(13414) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13414)))) severity failure;
    assert RAM(13415) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13415)))) severity failure;
    assert RAM(13416) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13416)))) severity failure;
    assert RAM(13417) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13417)))) severity failure;
    assert RAM(13418) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13418)))) severity failure;
    assert RAM(13419) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13419)))) severity failure;
    assert RAM(13420) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13420)))) severity failure;
    assert RAM(13421) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13421)))) severity failure;
    assert RAM(13422) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13422)))) severity failure;
    assert RAM(13423) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13423)))) severity failure;
    assert RAM(13424) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13424)))) severity failure;
    assert RAM(13425) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13425)))) severity failure;
    assert RAM(13426) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13426)))) severity failure;
    assert RAM(13427) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13427)))) severity failure;
    assert RAM(13428) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13428)))) severity failure;
    assert RAM(13429) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13429)))) severity failure;
    assert RAM(13430) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(13430)))) severity failure;
    assert RAM(13431) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13431)))) severity failure;
    assert RAM(13432) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13432)))) severity failure;
    assert RAM(13433) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(13433)))) severity failure;

    assert false report "Simulation Ended! TEST PASSATO" severity failure;
end process test;

end shlev7tb;
