-------------------------------------------------------------------------------
--
-- Final examination - Digital Logic Design
-- Alberto Boffi - Politecnico di Milano, AY 2020/21
-- TEST MODULE: Shift level = 4
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity shlev4_tb is
end shlev4_tb;

architecture shlev4tb of shlev4_tb is
constant c_CLOCK_PERIOD         : time := 15 ns;
signal   tb_done                : std_logic;
signal   mem_address            : std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst                 : std_logic := '0';
signal   tb_start               : std_logic := '0';
signal   tb_clk                 : std_logic := '0';
signal   mem_o_data,mem_i_data  : std_logic_vector (7 downto 0);
signal   enable_wire            : std_logic;
signal   mem_we                 : std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);


signal RAM: ram_type :=
	(0 => std_logic_vector(to_unsigned(111, 8)),
	1 => std_logic_vector(to_unsigned(8, 8)),
	2 => std_logic_vector(to_unsigned(150, 8)),
	3 => std_logic_vector(to_unsigned(163, 8)),
	4 => std_logic_vector(to_unsigned(159, 8)),
	5 => std_logic_vector(to_unsigned(155, 8)),
	6 => std_logic_vector(to_unsigned(159, 8)),
	7 => std_logic_vector(to_unsigned(154, 8)),
	8 => std_logic_vector(to_unsigned(159, 8)),
	9 => std_logic_vector(to_unsigned(152, 8)),
	10 => std_logic_vector(to_unsigned(155, 8)),
	11 => std_logic_vector(to_unsigned(162, 8)),
	12 => std_logic_vector(to_unsigned(157, 8)),
	13 => std_logic_vector(to_unsigned(166, 8)),
	14 => std_logic_vector(to_unsigned(159, 8)),
	15 => std_logic_vector(to_unsigned(165, 8)),
	16 => std_logic_vector(to_unsigned(150, 8)),
	17 => std_logic_vector(to_unsigned(154, 8)),
	18 => std_logic_vector(to_unsigned(159, 8)),
	19 => std_logic_vector(to_unsigned(159, 8)),
	20 => std_logic_vector(to_unsigned(154, 8)),
	21 => std_logic_vector(to_unsigned(155, 8)),
	22 => std_logic_vector(to_unsigned(165, 8)),
	23 => std_logic_vector(to_unsigned(157, 8)),
	24 => std_logic_vector(to_unsigned(160, 8)),
	25 => std_logic_vector(to_unsigned(153, 8)),
	26 => std_logic_vector(to_unsigned(164, 8)),
	27 => std_logic_vector(to_unsigned(163, 8)),
	28 => std_logic_vector(to_unsigned(160, 8)),
	29 => std_logic_vector(to_unsigned(158, 8)),
	30 => std_logic_vector(to_unsigned(151, 8)),
	31 => std_logic_vector(to_unsigned(160, 8)),
	32 => std_logic_vector(to_unsigned(162, 8)),
	33 => std_logic_vector(to_unsigned(160, 8)),
	34 => std_logic_vector(to_unsigned(165, 8)),
	35 => std_logic_vector(to_unsigned(163, 8)),
	36 => std_logic_vector(to_unsigned(152, 8)),
	37 => std_logic_vector(to_unsigned(149, 8)),
	38 => std_logic_vector(to_unsigned(160, 8)),
	39 => std_logic_vector(to_unsigned(158, 8)),
	40 => std_logic_vector(to_unsigned(149, 8)),
	41 => std_logic_vector(to_unsigned(152, 8)),
	42 => std_logic_vector(to_unsigned(149, 8)),
	43 => std_logic_vector(to_unsigned(153, 8)),
	44 => std_logic_vector(to_unsigned(153, 8)),
	45 => std_logic_vector(to_unsigned(159, 8)),
	46 => std_logic_vector(to_unsigned(152, 8)),
	47 => std_logic_vector(to_unsigned(152, 8)),
	48 => std_logic_vector(to_unsigned(161, 8)),
	49 => std_logic_vector(to_unsigned(155, 8)),
	50 => std_logic_vector(to_unsigned(156, 8)),
	51 => std_logic_vector(to_unsigned(150, 8)),
	52 => std_logic_vector(to_unsigned(160, 8)),
	53 => std_logic_vector(to_unsigned(155, 8)),
	54 => std_logic_vector(to_unsigned(163, 8)),
	55 => std_logic_vector(to_unsigned(161, 8)),
	56 => std_logic_vector(to_unsigned(164, 8)),
	57 => std_logic_vector(to_unsigned(165, 8)),
	58 => std_logic_vector(to_unsigned(150, 8)),
	59 => std_logic_vector(to_unsigned(159, 8)),
	60 => std_logic_vector(to_unsigned(155, 8)),
	61 => std_logic_vector(to_unsigned(166, 8)),
	62 => std_logic_vector(to_unsigned(155, 8)),
	63 => std_logic_vector(to_unsigned(159, 8)),
	64 => std_logic_vector(to_unsigned(162, 8)),
	65 => std_logic_vector(to_unsigned(163, 8)),
	66 => std_logic_vector(to_unsigned(151, 8)),
	67 => std_logic_vector(to_unsigned(160, 8)),
	68 => std_logic_vector(to_unsigned(163, 8)),
	69 => std_logic_vector(to_unsigned(159, 8)),
	70 => std_logic_vector(to_unsigned(165, 8)),
	71 => std_logic_vector(to_unsigned(151, 8)),
	72 => std_logic_vector(to_unsigned(159, 8)),
	73 => std_logic_vector(to_unsigned(152, 8)),
	74 => std_logic_vector(to_unsigned(165, 8)),
	75 => std_logic_vector(to_unsigned(153, 8)),
	76 => std_logic_vector(to_unsigned(160, 8)),
	77 => std_logic_vector(to_unsigned(157, 8)),
	78 => std_logic_vector(to_unsigned(153, 8)),
	79 => std_logic_vector(to_unsigned(165, 8)),
	80 => std_logic_vector(to_unsigned(151, 8)),
	81 => std_logic_vector(to_unsigned(152, 8)),
	82 => std_logic_vector(to_unsigned(162, 8)),
	83 => std_logic_vector(to_unsigned(162, 8)),
	84 => std_logic_vector(to_unsigned(161, 8)),
	85 => std_logic_vector(to_unsigned(160, 8)),
	86 => std_logic_vector(to_unsigned(165, 8)),
	87 => std_logic_vector(to_unsigned(155, 8)),
	88 => std_logic_vector(to_unsigned(164, 8)),
	89 => std_logic_vector(to_unsigned(149, 8)),
	90 => std_logic_vector(to_unsigned(166, 8)),
	91 => std_logic_vector(to_unsigned(164, 8)),
	92 => std_logic_vector(to_unsigned(156, 8)),
	93 => std_logic_vector(to_unsigned(159, 8)),
	94 => std_logic_vector(to_unsigned(152, 8)),
	95 => std_logic_vector(to_unsigned(156, 8)),
	96 => std_logic_vector(to_unsigned(158, 8)),
	97 => std_logic_vector(to_unsigned(150, 8)),
	98 => std_logic_vector(to_unsigned(150, 8)),
	99 => std_logic_vector(to_unsigned(162, 8)),
	100 => std_logic_vector(to_unsigned(151, 8)),
	101 => std_logic_vector(to_unsigned(157, 8)),
	102 => std_logic_vector(to_unsigned(159, 8)),
	103 => std_logic_vector(to_unsigned(149, 8)),
	104 => std_logic_vector(to_unsigned(165, 8)),
	105 => std_logic_vector(to_unsigned(150, 8)),
	106 => std_logic_vector(to_unsigned(163, 8)),
	107 => std_logic_vector(to_unsigned(155, 8)),
	108 => std_logic_vector(to_unsigned(150, 8)),
	109 => std_logic_vector(to_unsigned(161, 8)),
	110 => std_logic_vector(to_unsigned(162, 8)),
	111 => std_logic_vector(to_unsigned(155, 8)),
	112 => std_logic_vector(to_unsigned(163, 8)),
	113 => std_logic_vector(to_unsigned(161, 8)),
	114 => std_logic_vector(to_unsigned(163, 8)),
	115 => std_logic_vector(to_unsigned(156, 8)),
	116 => std_logic_vector(to_unsigned(156, 8)),
	117 => std_logic_vector(to_unsigned(151, 8)),
	118 => std_logic_vector(to_unsigned(151, 8)),
	119 => std_logic_vector(to_unsigned(154, 8)),
	120 => std_logic_vector(to_unsigned(164, 8)),
	121 => std_logic_vector(to_unsigned(153, 8)),
	122 => std_logic_vector(to_unsigned(158, 8)),
	123 => std_logic_vector(to_unsigned(166, 8)),
	124 => std_logic_vector(to_unsigned(155, 8)),
	125 => std_logic_vector(to_unsigned(160, 8)),
	126 => std_logic_vector(to_unsigned(155, 8)),
	127 => std_logic_vector(to_unsigned(160, 8)),
	128 => std_logic_vector(to_unsigned(156, 8)),
	129 => std_logic_vector(to_unsigned(164, 8)),
	130 => std_logic_vector(to_unsigned(153, 8)),
	131 => std_logic_vector(to_unsigned(158, 8)),
	132 => std_logic_vector(to_unsigned(159, 8)),
	133 => std_logic_vector(to_unsigned(157, 8)),
	134 => std_logic_vector(to_unsigned(162, 8)),
	135 => std_logic_vector(to_unsigned(164, 8)),
	136 => std_logic_vector(to_unsigned(164, 8)),
	137 => std_logic_vector(to_unsigned(149, 8)),
	138 => std_logic_vector(to_unsigned(158, 8)),
	139 => std_logic_vector(to_unsigned(156, 8)),
	140 => std_logic_vector(to_unsigned(166, 8)),
	141 => std_logic_vector(to_unsigned(155, 8)),
	142 => std_logic_vector(to_unsigned(160, 8)),
	143 => std_logic_vector(to_unsigned(158, 8)),
	144 => std_logic_vector(to_unsigned(151, 8)),
	145 => std_logic_vector(to_unsigned(152, 8)),
	146 => std_logic_vector(to_unsigned(162, 8)),
	147 => std_logic_vector(to_unsigned(162, 8)),
	148 => std_logic_vector(to_unsigned(153, 8)),
	149 => std_logic_vector(to_unsigned(149, 8)),
	150 => std_logic_vector(to_unsigned(153, 8)),
	151 => std_logic_vector(to_unsigned(149, 8)),
	152 => std_logic_vector(to_unsigned(152, 8)),
	153 => std_logic_vector(to_unsigned(152, 8)),
	154 => std_logic_vector(to_unsigned(155, 8)),
	155 => std_logic_vector(to_unsigned(159, 8)),
	156 => std_logic_vector(to_unsigned(158, 8)),
	157 => std_logic_vector(to_unsigned(159, 8)),
	158 => std_logic_vector(to_unsigned(165, 8)),
	159 => std_logic_vector(to_unsigned(151, 8)),
	160 => std_logic_vector(to_unsigned(150, 8)),
	161 => std_logic_vector(to_unsigned(153, 8)),
	162 => std_logic_vector(to_unsigned(166, 8)),
	163 => std_logic_vector(to_unsigned(152, 8)),
	164 => std_logic_vector(to_unsigned(150, 8)),
	165 => std_logic_vector(to_unsigned(155, 8)),
	166 => std_logic_vector(to_unsigned(159, 8)),
	167 => std_logic_vector(to_unsigned(150, 8)),
	168 => std_logic_vector(to_unsigned(155, 8)),
	169 => std_logic_vector(to_unsigned(152, 8)),
	170 => std_logic_vector(to_unsigned(150, 8)),
	171 => std_logic_vector(to_unsigned(151, 8)),
	172 => std_logic_vector(to_unsigned(163, 8)),
	173 => std_logic_vector(to_unsigned(155, 8)),
	174 => std_logic_vector(to_unsigned(164, 8)),
	175 => std_logic_vector(to_unsigned(151, 8)),
	176 => std_logic_vector(to_unsigned(164, 8)),
	177 => std_logic_vector(to_unsigned(157, 8)),
	178 => std_logic_vector(to_unsigned(157, 8)),
	179 => std_logic_vector(to_unsigned(164, 8)),
	180 => std_logic_vector(to_unsigned(166, 8)),
	181 => std_logic_vector(to_unsigned(160, 8)),
	182 => std_logic_vector(to_unsigned(150, 8)),
	183 => std_logic_vector(to_unsigned(162, 8)),
	184 => std_logic_vector(to_unsigned(160, 8)),
	185 => std_logic_vector(to_unsigned(165, 8)),
	186 => std_logic_vector(to_unsigned(150, 8)),
	187 => std_logic_vector(to_unsigned(157, 8)),
	188 => std_logic_vector(to_unsigned(151, 8)),
	189 => std_logic_vector(to_unsigned(152, 8)),
	190 => std_logic_vector(to_unsigned(154, 8)),
	191 => std_logic_vector(to_unsigned(153, 8)),
	192 => std_logic_vector(to_unsigned(152, 8)),
	193 => std_logic_vector(to_unsigned(149, 8)),
	194 => std_logic_vector(to_unsigned(151, 8)),
	195 => std_logic_vector(to_unsigned(162, 8)),
	196 => std_logic_vector(to_unsigned(152, 8)),
	197 => std_logic_vector(to_unsigned(150, 8)),
	198 => std_logic_vector(to_unsigned(163, 8)),
	199 => std_logic_vector(to_unsigned(160, 8)),
	200 => std_logic_vector(to_unsigned(165, 8)),
	201 => std_logic_vector(to_unsigned(151, 8)),
	202 => std_logic_vector(to_unsigned(165, 8)),
	203 => std_logic_vector(to_unsigned(152, 8)),
	204 => std_logic_vector(to_unsigned(150, 8)),
	205 => std_logic_vector(to_unsigned(150, 8)),
	206 => std_logic_vector(to_unsigned(152, 8)),
	207 => std_logic_vector(to_unsigned(157, 8)),
	208 => std_logic_vector(to_unsigned(154, 8)),
	209 => std_logic_vector(to_unsigned(151, 8)),
	210 => std_logic_vector(to_unsigned(164, 8)),
	211 => std_logic_vector(to_unsigned(149, 8)),
	212 => std_logic_vector(to_unsigned(153, 8)),
	213 => std_logic_vector(to_unsigned(166, 8)),
	214 => std_logic_vector(to_unsigned(149, 8)),
	215 => std_logic_vector(to_unsigned(152, 8)),
	216 => std_logic_vector(to_unsigned(165, 8)),
	217 => std_logic_vector(to_unsigned(152, 8)),
	218 => std_logic_vector(to_unsigned(156, 8)),
	219 => std_logic_vector(to_unsigned(160, 8)),
	220 => std_logic_vector(to_unsigned(165, 8)),
	221 => std_logic_vector(to_unsigned(150, 8)),
	222 => std_logic_vector(to_unsigned(154, 8)),
	223 => std_logic_vector(to_unsigned(152, 8)),
	224 => std_logic_vector(to_unsigned(164, 8)),
	225 => std_logic_vector(to_unsigned(150, 8)),
	226 => std_logic_vector(to_unsigned(165, 8)),
	227 => std_logic_vector(to_unsigned(159, 8)),
	228 => std_logic_vector(to_unsigned(162, 8)),
	229 => std_logic_vector(to_unsigned(158, 8)),
	230 => std_logic_vector(to_unsigned(166, 8)),
	231 => std_logic_vector(to_unsigned(165, 8)),
	232 => std_logic_vector(to_unsigned(155, 8)),
	233 => std_logic_vector(to_unsigned(155, 8)),
	234 => std_logic_vector(to_unsigned(158, 8)),
	235 => std_logic_vector(to_unsigned(166, 8)),
	236 => std_logic_vector(to_unsigned(154, 8)),
	237 => std_logic_vector(to_unsigned(153, 8)),
	238 => std_logic_vector(to_unsigned(154, 8)),
	239 => std_logic_vector(to_unsigned(157, 8)),
	240 => std_logic_vector(to_unsigned(160, 8)),
	241 => std_logic_vector(to_unsigned(160, 8)),
	242 => std_logic_vector(to_unsigned(152, 8)),
	243 => std_logic_vector(to_unsigned(166, 8)),
	244 => std_logic_vector(to_unsigned(164, 8)),
	245 => std_logic_vector(to_unsigned(165, 8)),
	246 => std_logic_vector(to_unsigned(161, 8)),
	247 => std_logic_vector(to_unsigned(156, 8)),
	248 => std_logic_vector(to_unsigned(152, 8)),
	249 => std_logic_vector(to_unsigned(160, 8)),
	250 => std_logic_vector(to_unsigned(163, 8)),
	251 => std_logic_vector(to_unsigned(150, 8)),
	252 => std_logic_vector(to_unsigned(166, 8)),
	253 => std_logic_vector(to_unsigned(150, 8)),
	254 => std_logic_vector(to_unsigned(149, 8)),
	255 => std_logic_vector(to_unsigned(150, 8)),
	256 => std_logic_vector(to_unsigned(165, 8)),
	257 => std_logic_vector(to_unsigned(166, 8)),
	258 => std_logic_vector(to_unsigned(166, 8)),
	259 => std_logic_vector(to_unsigned(149, 8)),
	260 => std_logic_vector(to_unsigned(164, 8)),
	261 => std_logic_vector(to_unsigned(160, 8)),
	262 => std_logic_vector(to_unsigned(153, 8)),
	263 => std_logic_vector(to_unsigned(166, 8)),
	264 => std_logic_vector(to_unsigned(159, 8)),
	265 => std_logic_vector(to_unsigned(158, 8)),
	266 => std_logic_vector(to_unsigned(158, 8)),
	267 => std_logic_vector(to_unsigned(149, 8)),
	268 => std_logic_vector(to_unsigned(166, 8)),
	269 => std_logic_vector(to_unsigned(151, 8)),
	270 => std_logic_vector(to_unsigned(158, 8)),
	271 => std_logic_vector(to_unsigned(156, 8)),
	272 => std_logic_vector(to_unsigned(153, 8)),
	273 => std_logic_vector(to_unsigned(165, 8)),
	274 => std_logic_vector(to_unsigned(156, 8)),
	275 => std_logic_vector(to_unsigned(165, 8)),
	276 => std_logic_vector(to_unsigned(162, 8)),
	277 => std_logic_vector(to_unsigned(157, 8)),
	278 => std_logic_vector(to_unsigned(154, 8)),
	279 => std_logic_vector(to_unsigned(162, 8)),
	280 => std_logic_vector(to_unsigned(159, 8)),
	281 => std_logic_vector(to_unsigned(160, 8)),
	282 => std_logic_vector(to_unsigned(151, 8)),
	283 => std_logic_vector(to_unsigned(157, 8)),
	284 => std_logic_vector(to_unsigned(157, 8)),
	285 => std_logic_vector(to_unsigned(153, 8)),
	286 => std_logic_vector(to_unsigned(155, 8)),
	287 => std_logic_vector(to_unsigned(159, 8)),
	288 => std_logic_vector(to_unsigned(162, 8)),
	289 => std_logic_vector(to_unsigned(163, 8)),
	290 => std_logic_vector(to_unsigned(150, 8)),
	291 => std_logic_vector(to_unsigned(166, 8)),
	292 => std_logic_vector(to_unsigned(166, 8)),
	293 => std_logic_vector(to_unsigned(165, 8)),
	294 => std_logic_vector(to_unsigned(154, 8)),
	295 => std_logic_vector(to_unsigned(153, 8)),
	296 => std_logic_vector(to_unsigned(157, 8)),
	297 => std_logic_vector(to_unsigned(152, 8)),
	298 => std_logic_vector(to_unsigned(166, 8)),
	299 => std_logic_vector(to_unsigned(151, 8)),
	300 => std_logic_vector(to_unsigned(153, 8)),
	301 => std_logic_vector(to_unsigned(162, 8)),
	302 => std_logic_vector(to_unsigned(151, 8)),
	303 => std_logic_vector(to_unsigned(149, 8)),
	304 => std_logic_vector(to_unsigned(160, 8)),
	305 => std_logic_vector(to_unsigned(161, 8)),
	306 => std_logic_vector(to_unsigned(151, 8)),
	307 => std_logic_vector(to_unsigned(149, 8)),
	308 => std_logic_vector(to_unsigned(162, 8)),
	309 => std_logic_vector(to_unsigned(163, 8)),
	310 => std_logic_vector(to_unsigned(163, 8)),
	311 => std_logic_vector(to_unsigned(150, 8)),
	312 => std_logic_vector(to_unsigned(160, 8)),
	313 => std_logic_vector(to_unsigned(153, 8)),
	314 => std_logic_vector(to_unsigned(159, 8)),
	315 => std_logic_vector(to_unsigned(166, 8)),
	316 => std_logic_vector(to_unsigned(162, 8)),
	317 => std_logic_vector(to_unsigned(150, 8)),
	318 => std_logic_vector(to_unsigned(150, 8)),
	319 => std_logic_vector(to_unsigned(153, 8)),
	320 => std_logic_vector(to_unsigned(156, 8)),
	321 => std_logic_vector(to_unsigned(162, 8)),
	322 => std_logic_vector(to_unsigned(158, 8)),
	323 => std_logic_vector(to_unsigned(164, 8)),
	324 => std_logic_vector(to_unsigned(149, 8)),
	325 => std_logic_vector(to_unsigned(149, 8)),
	326 => std_logic_vector(to_unsigned(151, 8)),
	327 => std_logic_vector(to_unsigned(155, 8)),
	328 => std_logic_vector(to_unsigned(159, 8)),
	329 => std_logic_vector(to_unsigned(153, 8)),
	330 => std_logic_vector(to_unsigned(158, 8)),
	331 => std_logic_vector(to_unsigned(160, 8)),
	332 => std_logic_vector(to_unsigned(154, 8)),
	333 => std_logic_vector(to_unsigned(164, 8)),
	334 => std_logic_vector(to_unsigned(152, 8)),
	335 => std_logic_vector(to_unsigned(153, 8)),
	336 => std_logic_vector(to_unsigned(150, 8)),
	337 => std_logic_vector(to_unsigned(163, 8)),
	338 => std_logic_vector(to_unsigned(164, 8)),
	339 => std_logic_vector(to_unsigned(153, 8)),
	340 => std_logic_vector(to_unsigned(166, 8)),
	341 => std_logic_vector(to_unsigned(151, 8)),
	342 => std_logic_vector(to_unsigned(155, 8)),
	343 => std_logic_vector(to_unsigned(152, 8)),
	344 => std_logic_vector(to_unsigned(163, 8)),
	345 => std_logic_vector(to_unsigned(161, 8)),
	346 => std_logic_vector(to_unsigned(160, 8)),
	347 => std_logic_vector(to_unsigned(164, 8)),
	348 => std_logic_vector(to_unsigned(154, 8)),
	349 => std_logic_vector(to_unsigned(161, 8)),
	350 => std_logic_vector(to_unsigned(161, 8)),
	351 => std_logic_vector(to_unsigned(165, 8)),
	352 => std_logic_vector(to_unsigned(161, 8)),
	353 => std_logic_vector(to_unsigned(157, 8)),
	354 => std_logic_vector(to_unsigned(161, 8)),
	355 => std_logic_vector(to_unsigned(156, 8)),
	356 => std_logic_vector(to_unsigned(162, 8)),
	357 => std_logic_vector(to_unsigned(156, 8)),
	358 => std_logic_vector(to_unsigned(165, 8)),
	359 => std_logic_vector(to_unsigned(158, 8)),
	360 => std_logic_vector(to_unsigned(149, 8)),
	361 => std_logic_vector(to_unsigned(164, 8)),
	362 => std_logic_vector(to_unsigned(152, 8)),
	363 => std_logic_vector(to_unsigned(150, 8)),
	364 => std_logic_vector(to_unsigned(165, 8)),
	365 => std_logic_vector(to_unsigned(155, 8)),
	366 => std_logic_vector(to_unsigned(156, 8)),
	367 => std_logic_vector(to_unsigned(153, 8)),
	368 => std_logic_vector(to_unsigned(160, 8)),
	369 => std_logic_vector(to_unsigned(155, 8)),
	370 => std_logic_vector(to_unsigned(154, 8)),
	371 => std_logic_vector(to_unsigned(152, 8)),
	372 => std_logic_vector(to_unsigned(160, 8)),
	373 => std_logic_vector(to_unsigned(163, 8)),
	374 => std_logic_vector(to_unsigned(165, 8)),
	375 => std_logic_vector(to_unsigned(159, 8)),
	376 => std_logic_vector(to_unsigned(166, 8)),
	377 => std_logic_vector(to_unsigned(161, 8)),
	378 => std_logic_vector(to_unsigned(157, 8)),
	379 => std_logic_vector(to_unsigned(156, 8)),
	380 => std_logic_vector(to_unsigned(162, 8)),
	381 => std_logic_vector(to_unsigned(154, 8)),
	382 => std_logic_vector(to_unsigned(159, 8)),
	383 => std_logic_vector(to_unsigned(156, 8)),
	384 => std_logic_vector(to_unsigned(149, 8)),
	385 => std_logic_vector(to_unsigned(158, 8)),
	386 => std_logic_vector(to_unsigned(166, 8)),
	387 => std_logic_vector(to_unsigned(157, 8)),
	388 => std_logic_vector(to_unsigned(156, 8)),
	389 => std_logic_vector(to_unsigned(153, 8)),
	390 => std_logic_vector(to_unsigned(150, 8)),
	391 => std_logic_vector(to_unsigned(157, 8)),
	392 => std_logic_vector(to_unsigned(156, 8)),
	393 => std_logic_vector(to_unsigned(159, 8)),
	394 => std_logic_vector(to_unsigned(151, 8)),
	395 => std_logic_vector(to_unsigned(149, 8)),
	396 => std_logic_vector(to_unsigned(151, 8)),
	397 => std_logic_vector(to_unsigned(164, 8)),
	398 => std_logic_vector(to_unsigned(165, 8)),
	399 => std_logic_vector(to_unsigned(151, 8)),
	400 => std_logic_vector(to_unsigned(161, 8)),
	401 => std_logic_vector(to_unsigned(161, 8)),
	402 => std_logic_vector(to_unsigned(154, 8)),
	403 => std_logic_vector(to_unsigned(155, 8)),
	404 => std_logic_vector(to_unsigned(165, 8)),
	405 => std_logic_vector(to_unsigned(155, 8)),
	406 => std_logic_vector(to_unsigned(161, 8)),
	407 => std_logic_vector(to_unsigned(155, 8)),
	408 => std_logic_vector(to_unsigned(165, 8)),
	409 => std_logic_vector(to_unsigned(160, 8)),
	410 => std_logic_vector(to_unsigned(159, 8)),
	411 => std_logic_vector(to_unsigned(159, 8)),
	412 => std_logic_vector(to_unsigned(159, 8)),
	413 => std_logic_vector(to_unsigned(162, 8)),
	414 => std_logic_vector(to_unsigned(151, 8)),
	415 => std_logic_vector(to_unsigned(158, 8)),
	416 => std_logic_vector(to_unsigned(165, 8)),
	417 => std_logic_vector(to_unsigned(166, 8)),
	418 => std_logic_vector(to_unsigned(165, 8)),
	419 => std_logic_vector(to_unsigned(154, 8)),
	420 => std_logic_vector(to_unsigned(158, 8)),
	421 => std_logic_vector(to_unsigned(153, 8)),
	422 => std_logic_vector(to_unsigned(160, 8)),
	423 => std_logic_vector(to_unsigned(152, 8)),
	424 => std_logic_vector(to_unsigned(160, 8)),
	425 => std_logic_vector(to_unsigned(159, 8)),
	426 => std_logic_vector(to_unsigned(154, 8)),
	427 => std_logic_vector(to_unsigned(162, 8)),
	428 => std_logic_vector(to_unsigned(153, 8)),
	429 => std_logic_vector(to_unsigned(166, 8)),
	430 => std_logic_vector(to_unsigned(155, 8)),
	431 => std_logic_vector(to_unsigned(152, 8)),
	432 => std_logic_vector(to_unsigned(162, 8)),
	433 => std_logic_vector(to_unsigned(153, 8)),
	434 => std_logic_vector(to_unsigned(161, 8)),
	435 => std_logic_vector(to_unsigned(159, 8)),
	436 => std_logic_vector(to_unsigned(155, 8)),
	437 => std_logic_vector(to_unsigned(157, 8)),
	438 => std_logic_vector(to_unsigned(151, 8)),
	439 => std_logic_vector(to_unsigned(164, 8)),
	440 => std_logic_vector(to_unsigned(152, 8)),
	441 => std_logic_vector(to_unsigned(150, 8)),
	442 => std_logic_vector(to_unsigned(160, 8)),
	443 => std_logic_vector(to_unsigned(163, 8)),
	444 => std_logic_vector(to_unsigned(152, 8)),
	445 => std_logic_vector(to_unsigned(151, 8)),
	446 => std_logic_vector(to_unsigned(154, 8)),
	447 => std_logic_vector(to_unsigned(149, 8)),
	448 => std_logic_vector(to_unsigned(158, 8)),
	449 => std_logic_vector(to_unsigned(163, 8)),
	450 => std_logic_vector(to_unsigned(151, 8)),
	451 => std_logic_vector(to_unsigned(149, 8)),
	452 => std_logic_vector(to_unsigned(164, 8)),
	453 => std_logic_vector(to_unsigned(156, 8)),
	454 => std_logic_vector(to_unsigned(160, 8)),
	455 => std_logic_vector(to_unsigned(159, 8)),
	456 => std_logic_vector(to_unsigned(166, 8)),
	457 => std_logic_vector(to_unsigned(151, 8)),
	458 => std_logic_vector(to_unsigned(165, 8)),
	459 => std_logic_vector(to_unsigned(162, 8)),
	460 => std_logic_vector(to_unsigned(158, 8)),
	461 => std_logic_vector(to_unsigned(161, 8)),
	462 => std_logic_vector(to_unsigned(151, 8)),
	463 => std_logic_vector(to_unsigned(161, 8)),
	464 => std_logic_vector(to_unsigned(161, 8)),
	465 => std_logic_vector(to_unsigned(154, 8)),
	466 => std_logic_vector(to_unsigned(150, 8)),
	467 => std_logic_vector(to_unsigned(165, 8)),
	468 => std_logic_vector(to_unsigned(154, 8)),
	469 => std_logic_vector(to_unsigned(153, 8)),
	470 => std_logic_vector(to_unsigned(165, 8)),
	471 => std_logic_vector(to_unsigned(164, 8)),
	472 => std_logic_vector(to_unsigned(150, 8)),
	473 => std_logic_vector(to_unsigned(160, 8)),
	474 => std_logic_vector(to_unsigned(163, 8)),
	475 => std_logic_vector(to_unsigned(153, 8)),
	476 => std_logic_vector(to_unsigned(163, 8)),
	477 => std_logic_vector(to_unsigned(166, 8)),
	478 => std_logic_vector(to_unsigned(151, 8)),
	479 => std_logic_vector(to_unsigned(158, 8)),
	480 => std_logic_vector(to_unsigned(154, 8)),
	481 => std_logic_vector(to_unsigned(158, 8)),
	482 => std_logic_vector(to_unsigned(161, 8)),
	483 => std_logic_vector(to_unsigned(164, 8)),
	484 => std_logic_vector(to_unsigned(154, 8)),
	485 => std_logic_vector(to_unsigned(151, 8)),
	486 => std_logic_vector(to_unsigned(158, 8)),
	487 => std_logic_vector(to_unsigned(158, 8)),
	488 => std_logic_vector(to_unsigned(162, 8)),
	489 => std_logic_vector(to_unsigned(160, 8)),
	490 => std_logic_vector(to_unsigned(155, 8)),
	491 => std_logic_vector(to_unsigned(161, 8)),
	492 => std_logic_vector(to_unsigned(152, 8)),
	493 => std_logic_vector(to_unsigned(161, 8)),
	494 => std_logic_vector(to_unsigned(154, 8)),
	495 => std_logic_vector(to_unsigned(164, 8)),
	496 => std_logic_vector(to_unsigned(166, 8)),
	497 => std_logic_vector(to_unsigned(159, 8)),
	498 => std_logic_vector(to_unsigned(160, 8)),
	499 => std_logic_vector(to_unsigned(154, 8)),
	500 => std_logic_vector(to_unsigned(163, 8)),
	501 => std_logic_vector(to_unsigned(149, 8)),
	502 => std_logic_vector(to_unsigned(166, 8)),
	503 => std_logic_vector(to_unsigned(166, 8)),
	504 => std_logic_vector(to_unsigned(157, 8)),
	505 => std_logic_vector(to_unsigned(152, 8)),
	506 => std_logic_vector(to_unsigned(159, 8)),
	507 => std_logic_vector(to_unsigned(158, 8)),
	508 => std_logic_vector(to_unsigned(163, 8)),
	509 => std_logic_vector(to_unsigned(155, 8)),
	510 => std_logic_vector(to_unsigned(156, 8)),
	511 => std_logic_vector(to_unsigned(153, 8)),
	512 => std_logic_vector(to_unsigned(165, 8)),
	513 => std_logic_vector(to_unsigned(162, 8)),
	514 => std_logic_vector(to_unsigned(153, 8)),
	515 => std_logic_vector(to_unsigned(161, 8)),
	516 => std_logic_vector(to_unsigned(164, 8)),
	517 => std_logic_vector(to_unsigned(150, 8)),
	518 => std_logic_vector(to_unsigned(163, 8)),
	519 => std_logic_vector(to_unsigned(165, 8)),
	520 => std_logic_vector(to_unsigned(163, 8)),
	521 => std_logic_vector(to_unsigned(161, 8)),
	522 => std_logic_vector(to_unsigned(162, 8)),
	523 => std_logic_vector(to_unsigned(165, 8)),
	524 => std_logic_vector(to_unsigned(158, 8)),
	525 => std_logic_vector(to_unsigned(152, 8)),
	526 => std_logic_vector(to_unsigned(152, 8)),
	527 => std_logic_vector(to_unsigned(165, 8)),
	528 => std_logic_vector(to_unsigned(163, 8)),
	529 => std_logic_vector(to_unsigned(157, 8)),
	530 => std_logic_vector(to_unsigned(153, 8)),
	531 => std_logic_vector(to_unsigned(160, 8)),
	532 => std_logic_vector(to_unsigned(161, 8)),
	533 => std_logic_vector(to_unsigned(159, 8)),
	534 => std_logic_vector(to_unsigned(157, 8)),
	535 => std_logic_vector(to_unsigned(152, 8)),
	536 => std_logic_vector(to_unsigned(158, 8)),
	537 => std_logic_vector(to_unsigned(156, 8)),
	538 => std_logic_vector(to_unsigned(161, 8)),
	539 => std_logic_vector(to_unsigned(160, 8)),
	540 => std_logic_vector(to_unsigned(158, 8)),
	541 => std_logic_vector(to_unsigned(151, 8)),
	542 => std_logic_vector(to_unsigned(150, 8)),
	543 => std_logic_vector(to_unsigned(152, 8)),
	544 => std_logic_vector(to_unsigned(151, 8)),
	545 => std_logic_vector(to_unsigned(150, 8)),
	546 => std_logic_vector(to_unsigned(154, 8)),
	547 => std_logic_vector(to_unsigned(165, 8)),
	548 => std_logic_vector(to_unsigned(160, 8)),
	549 => std_logic_vector(to_unsigned(150, 8)),
	550 => std_logic_vector(to_unsigned(161, 8)),
	551 => std_logic_vector(to_unsigned(153, 8)),
	552 => std_logic_vector(to_unsigned(158, 8)),
	553 => std_logic_vector(to_unsigned(152, 8)),
	554 => std_logic_vector(to_unsigned(159, 8)),
	555 => std_logic_vector(to_unsigned(156, 8)),
	556 => std_logic_vector(to_unsigned(161, 8)),
	557 => std_logic_vector(to_unsigned(157, 8)),
	558 => std_logic_vector(to_unsigned(150, 8)),
	559 => std_logic_vector(to_unsigned(151, 8)),
	560 => std_logic_vector(to_unsigned(163, 8)),
	561 => std_logic_vector(to_unsigned(152, 8)),
	562 => std_logic_vector(to_unsigned(154, 8)),
	563 => std_logic_vector(to_unsigned(163, 8)),
	564 => std_logic_vector(to_unsigned(160, 8)),
	565 => std_logic_vector(to_unsigned(152, 8)),
	566 => std_logic_vector(to_unsigned(154, 8)),
	567 => std_logic_vector(to_unsigned(159, 8)),
	568 => std_logic_vector(to_unsigned(160, 8)),
	569 => std_logic_vector(to_unsigned(166, 8)),
	570 => std_logic_vector(to_unsigned(161, 8)),
	571 => std_logic_vector(to_unsigned(164, 8)),
	572 => std_logic_vector(to_unsigned(160, 8)),
	573 => std_logic_vector(to_unsigned(164, 8)),
	574 => std_logic_vector(to_unsigned(165, 8)),
	575 => std_logic_vector(to_unsigned(166, 8)),
	576 => std_logic_vector(to_unsigned(152, 8)),
	577 => std_logic_vector(to_unsigned(158, 8)),
	578 => std_logic_vector(to_unsigned(164, 8)),
	579 => std_logic_vector(to_unsigned(165, 8)),
	580 => std_logic_vector(to_unsigned(155, 8)),
	581 => std_logic_vector(to_unsigned(157, 8)),
	582 => std_logic_vector(to_unsigned(159, 8)),
	583 => std_logic_vector(to_unsigned(151, 8)),
	584 => std_logic_vector(to_unsigned(158, 8)),
	585 => std_logic_vector(to_unsigned(152, 8)),
	586 => std_logic_vector(to_unsigned(165, 8)),
	587 => std_logic_vector(to_unsigned(153, 8)),
	588 => std_logic_vector(to_unsigned(151, 8)),
	589 => std_logic_vector(to_unsigned(156, 8)),
	590 => std_logic_vector(to_unsigned(161, 8)),
	591 => std_logic_vector(to_unsigned(154, 8)),
	592 => std_logic_vector(to_unsigned(163, 8)),
	593 => std_logic_vector(to_unsigned(160, 8)),
	594 => std_logic_vector(to_unsigned(150, 8)),
	595 => std_logic_vector(to_unsigned(149, 8)),
	596 => std_logic_vector(to_unsigned(166, 8)),
	597 => std_logic_vector(to_unsigned(151, 8)),
	598 => std_logic_vector(to_unsigned(155, 8)),
	599 => std_logic_vector(to_unsigned(166, 8)),
	600 => std_logic_vector(to_unsigned(164, 8)),
	601 => std_logic_vector(to_unsigned(161, 8)),
	602 => std_logic_vector(to_unsigned(157, 8)),
	603 => std_logic_vector(to_unsigned(153, 8)),
	604 => std_logic_vector(to_unsigned(157, 8)),
	605 => std_logic_vector(to_unsigned(162, 8)),
	606 => std_logic_vector(to_unsigned(162, 8)),
	607 => std_logic_vector(to_unsigned(165, 8)),
	608 => std_logic_vector(to_unsigned(151, 8)),
	609 => std_logic_vector(to_unsigned(152, 8)),
	610 => std_logic_vector(to_unsigned(152, 8)),
	611 => std_logic_vector(to_unsigned(156, 8)),
	612 => std_logic_vector(to_unsigned(155, 8)),
	613 => std_logic_vector(to_unsigned(153, 8)),
	614 => std_logic_vector(to_unsigned(154, 8)),
	615 => std_logic_vector(to_unsigned(155, 8)),
	616 => std_logic_vector(to_unsigned(161, 8)),
	617 => std_logic_vector(to_unsigned(165, 8)),
	618 => std_logic_vector(to_unsigned(150, 8)),
	619 => std_logic_vector(to_unsigned(156, 8)),
	620 => std_logic_vector(to_unsigned(166, 8)),
	621 => std_logic_vector(to_unsigned(156, 8)),
	622 => std_logic_vector(to_unsigned(156, 8)),
	623 => std_logic_vector(to_unsigned(165, 8)),
	624 => std_logic_vector(to_unsigned(155, 8)),
	625 => std_logic_vector(to_unsigned(162, 8)),
	626 => std_logic_vector(to_unsigned(151, 8)),
	627 => std_logic_vector(to_unsigned(164, 8)),
	628 => std_logic_vector(to_unsigned(158, 8)),
	629 => std_logic_vector(to_unsigned(159, 8)),
	630 => std_logic_vector(to_unsigned(163, 8)),
	631 => std_logic_vector(to_unsigned(161, 8)),
	632 => std_logic_vector(to_unsigned(160, 8)),
	633 => std_logic_vector(to_unsigned(163, 8)),
	634 => std_logic_vector(to_unsigned(161, 8)),
	635 => std_logic_vector(to_unsigned(153, 8)),
	636 => std_logic_vector(to_unsigned(158, 8)),
	637 => std_logic_vector(to_unsigned(153, 8)),
	638 => std_logic_vector(to_unsigned(163, 8)),
	639 => std_logic_vector(to_unsigned(152, 8)),
	640 => std_logic_vector(to_unsigned(152, 8)),
	641 => std_logic_vector(to_unsigned(153, 8)),
	642 => std_logic_vector(to_unsigned(160, 8)),
	643 => std_logic_vector(to_unsigned(157, 8)),
	644 => std_logic_vector(to_unsigned(150, 8)),
	645 => std_logic_vector(to_unsigned(164, 8)),
	646 => std_logic_vector(to_unsigned(164, 8)),
	647 => std_logic_vector(to_unsigned(155, 8)),
	648 => std_logic_vector(to_unsigned(160, 8)),
	649 => std_logic_vector(to_unsigned(165, 8)),
	650 => std_logic_vector(to_unsigned(157, 8)),
	651 => std_logic_vector(to_unsigned(149, 8)),
	652 => std_logic_vector(to_unsigned(162, 8)),
	653 => std_logic_vector(to_unsigned(165, 8)),
	654 => std_logic_vector(to_unsigned(157, 8)),
	655 => std_logic_vector(to_unsigned(165, 8)),
	656 => std_logic_vector(to_unsigned(150, 8)),
	657 => std_logic_vector(to_unsigned(158, 8)),
	658 => std_logic_vector(to_unsigned(163, 8)),
	659 => std_logic_vector(to_unsigned(157, 8)),
	660 => std_logic_vector(to_unsigned(161, 8)),
	661 => std_logic_vector(to_unsigned(162, 8)),
	662 => std_logic_vector(to_unsigned(160, 8)),
	663 => std_logic_vector(to_unsigned(159, 8)),
	664 => std_logic_vector(to_unsigned(149, 8)),
	665 => std_logic_vector(to_unsigned(166, 8)),
	666 => std_logic_vector(to_unsigned(159, 8)),
	667 => std_logic_vector(to_unsigned(150, 8)),
	668 => std_logic_vector(to_unsigned(155, 8)),
	669 => std_logic_vector(to_unsigned(166, 8)),
	670 => std_logic_vector(to_unsigned(157, 8)),
	671 => std_logic_vector(to_unsigned(158, 8)),
	672 => std_logic_vector(to_unsigned(156, 8)),
	673 => std_logic_vector(to_unsigned(163, 8)),
	674 => std_logic_vector(to_unsigned(157, 8)),
	675 => std_logic_vector(to_unsigned(157, 8)),
	676 => std_logic_vector(to_unsigned(166, 8)),
	677 => std_logic_vector(to_unsigned(158, 8)),
	678 => std_logic_vector(to_unsigned(150, 8)),
	679 => std_logic_vector(to_unsigned(150, 8)),
	680 => std_logic_vector(to_unsigned(159, 8)),
	681 => std_logic_vector(to_unsigned(151, 8)),
	682 => std_logic_vector(to_unsigned(164, 8)),
	683 => std_logic_vector(to_unsigned(160, 8)),
	684 => std_logic_vector(to_unsigned(151, 8)),
	685 => std_logic_vector(to_unsigned(164, 8)),
	686 => std_logic_vector(to_unsigned(163, 8)),
	687 => std_logic_vector(to_unsigned(157, 8)),
	688 => std_logic_vector(to_unsigned(165, 8)),
	689 => std_logic_vector(to_unsigned(150, 8)),
	690 => std_logic_vector(to_unsigned(160, 8)),
	691 => std_logic_vector(to_unsigned(159, 8)),
	692 => std_logic_vector(to_unsigned(163, 8)),
	693 => std_logic_vector(to_unsigned(149, 8)),
	694 => std_logic_vector(to_unsigned(162, 8)),
	695 => std_logic_vector(to_unsigned(157, 8)),
	696 => std_logic_vector(to_unsigned(166, 8)),
	697 => std_logic_vector(to_unsigned(158, 8)),
	698 => std_logic_vector(to_unsigned(155, 8)),
	699 => std_logic_vector(to_unsigned(150, 8)),
	700 => std_logic_vector(to_unsigned(165, 8)),
	701 => std_logic_vector(to_unsigned(150, 8)),
	702 => std_logic_vector(to_unsigned(161, 8)),
	703 => std_logic_vector(to_unsigned(165, 8)),
	704 => std_logic_vector(to_unsigned(162, 8)),
	705 => std_logic_vector(to_unsigned(165, 8)),
	706 => std_logic_vector(to_unsigned(150, 8)),
	707 => std_logic_vector(to_unsigned(155, 8)),
	708 => std_logic_vector(to_unsigned(162, 8)),
	709 => std_logic_vector(to_unsigned(162, 8)),
	710 => std_logic_vector(to_unsigned(152, 8)),
	711 => std_logic_vector(to_unsigned(155, 8)),
	712 => std_logic_vector(to_unsigned(165, 8)),
	713 => std_logic_vector(to_unsigned(161, 8)),
	714 => std_logic_vector(to_unsigned(157, 8)),
	715 => std_logic_vector(to_unsigned(157, 8)),
	716 => std_logic_vector(to_unsigned(159, 8)),
	717 => std_logic_vector(to_unsigned(153, 8)),
	718 => std_logic_vector(to_unsigned(154, 8)),
	719 => std_logic_vector(to_unsigned(159, 8)),
	720 => std_logic_vector(to_unsigned(163, 8)),
	721 => std_logic_vector(to_unsigned(154, 8)),
	722 => std_logic_vector(to_unsigned(165, 8)),
	723 => std_logic_vector(to_unsigned(163, 8)),
	724 => std_logic_vector(to_unsigned(153, 8)),
	725 => std_logic_vector(to_unsigned(159, 8)),
	726 => std_logic_vector(to_unsigned(155, 8)),
	727 => std_logic_vector(to_unsigned(154, 8)),
	728 => std_logic_vector(to_unsigned(150, 8)),
	729 => std_logic_vector(to_unsigned(161, 8)),
	730 => std_logic_vector(to_unsigned(152, 8)),
	731 => std_logic_vector(to_unsigned(158, 8)),
	732 => std_logic_vector(to_unsigned(158, 8)),
	733 => std_logic_vector(to_unsigned(162, 8)),
	734 => std_logic_vector(to_unsigned(164, 8)),
	735 => std_logic_vector(to_unsigned(151, 8)),
	736 => std_logic_vector(to_unsigned(153, 8)),
	737 => std_logic_vector(to_unsigned(156, 8)),
	738 => std_logic_vector(to_unsigned(163, 8)),
	739 => std_logic_vector(to_unsigned(162, 8)),
	740 => std_logic_vector(to_unsigned(149, 8)),
	741 => std_logic_vector(to_unsigned(165, 8)),
	742 => std_logic_vector(to_unsigned(160, 8)),
	743 => std_logic_vector(to_unsigned(155, 8)),
	744 => std_logic_vector(to_unsigned(162, 8)),
	745 => std_logic_vector(to_unsigned(159, 8)),
	746 => std_logic_vector(to_unsigned(154, 8)),
	747 => std_logic_vector(to_unsigned(155, 8)),
	748 => std_logic_vector(to_unsigned(150, 8)),
	749 => std_logic_vector(to_unsigned(162, 8)),
	750 => std_logic_vector(to_unsigned(152, 8)),
	751 => std_logic_vector(to_unsigned(164, 8)),
	752 => std_logic_vector(to_unsigned(165, 8)),
	753 => std_logic_vector(to_unsigned(165, 8)),
	754 => std_logic_vector(to_unsigned(155, 8)),
	755 => std_logic_vector(to_unsigned(153, 8)),
	756 => std_logic_vector(to_unsigned(165, 8)),
	757 => std_logic_vector(to_unsigned(159, 8)),
	758 => std_logic_vector(to_unsigned(166, 8)),
	759 => std_logic_vector(to_unsigned(158, 8)),
	760 => std_logic_vector(to_unsigned(156, 8)),
	761 => std_logic_vector(to_unsigned(151, 8)),
	762 => std_logic_vector(to_unsigned(159, 8)),
	763 => std_logic_vector(to_unsigned(149, 8)),
	764 => std_logic_vector(to_unsigned(158, 8)),
	765 => std_logic_vector(to_unsigned(159, 8)),
	766 => std_logic_vector(to_unsigned(152, 8)),
	767 => std_logic_vector(to_unsigned(157, 8)),
	768 => std_logic_vector(to_unsigned(160, 8)),
	769 => std_logic_vector(to_unsigned(159, 8)),
	770 => std_logic_vector(to_unsigned(155, 8)),
	771 => std_logic_vector(to_unsigned(150, 8)),
	772 => std_logic_vector(to_unsigned(166, 8)),
	773 => std_logic_vector(to_unsigned(163, 8)),
	774 => std_logic_vector(to_unsigned(161, 8)),
	775 => std_logic_vector(to_unsigned(159, 8)),
	776 => std_logic_vector(to_unsigned(160, 8)),
	777 => std_logic_vector(to_unsigned(150, 8)),
	778 => std_logic_vector(to_unsigned(154, 8)),
	779 => std_logic_vector(to_unsigned(164, 8)),
	780 => std_logic_vector(to_unsigned(151, 8)),
	781 => std_logic_vector(to_unsigned(159, 8)),
	782 => std_logic_vector(to_unsigned(154, 8)),
	783 => std_logic_vector(to_unsigned(153, 8)),
	784 => std_logic_vector(to_unsigned(154, 8)),
	785 => std_logic_vector(to_unsigned(165, 8)),
	786 => std_logic_vector(to_unsigned(159, 8)),
	787 => std_logic_vector(to_unsigned(159, 8)),
	788 => std_logic_vector(to_unsigned(162, 8)),
	789 => std_logic_vector(to_unsigned(151, 8)),
	790 => std_logic_vector(to_unsigned(164, 8)),
	791 => std_logic_vector(to_unsigned(150, 8)),
	792 => std_logic_vector(to_unsigned(160, 8)),
	793 => std_logic_vector(to_unsigned(161, 8)),
	794 => std_logic_vector(to_unsigned(164, 8)),
	795 => std_logic_vector(to_unsigned(164, 8)),
	796 => std_logic_vector(to_unsigned(157, 8)),
	797 => std_logic_vector(to_unsigned(153, 8)),
	798 => std_logic_vector(to_unsigned(159, 8)),
	799 => std_logic_vector(to_unsigned(165, 8)),
	800 => std_logic_vector(to_unsigned(158, 8)),
	801 => std_logic_vector(to_unsigned(153, 8)),
	802 => std_logic_vector(to_unsigned(151, 8)),
	803 => std_logic_vector(to_unsigned(150, 8)),
	804 => std_logic_vector(to_unsigned(157, 8)),
	805 => std_logic_vector(to_unsigned(150, 8)),
	806 => std_logic_vector(to_unsigned(149, 8)),
	807 => std_logic_vector(to_unsigned(159, 8)),
	808 => std_logic_vector(to_unsigned(161, 8)),
	809 => std_logic_vector(to_unsigned(159, 8)),
	810 => std_logic_vector(to_unsigned(162, 8)),
	811 => std_logic_vector(to_unsigned(164, 8)),
	812 => std_logic_vector(to_unsigned(157, 8)),
	813 => std_logic_vector(to_unsigned(165, 8)),
	814 => std_logic_vector(to_unsigned(160, 8)),
	815 => std_logic_vector(to_unsigned(153, 8)),
	816 => std_logic_vector(to_unsigned(161, 8)),
	817 => std_logic_vector(to_unsigned(162, 8)),
	818 => std_logic_vector(to_unsigned(166, 8)),
	819 => std_logic_vector(to_unsigned(166, 8)),
	820 => std_logic_vector(to_unsigned(152, 8)),
	821 => std_logic_vector(to_unsigned(151, 8)),
	822 => std_logic_vector(to_unsigned(160, 8)),
	823 => std_logic_vector(to_unsigned(159, 8)),
	824 => std_logic_vector(to_unsigned(151, 8)),
	825 => std_logic_vector(to_unsigned(158, 8)),
	826 => std_logic_vector(to_unsigned(149, 8)),
	827 => std_logic_vector(to_unsigned(151, 8)),
	828 => std_logic_vector(to_unsigned(159, 8)),
	829 => std_logic_vector(to_unsigned(151, 8)),
	830 => std_logic_vector(to_unsigned(164, 8)),
	831 => std_logic_vector(to_unsigned(162, 8)),
	832 => std_logic_vector(to_unsigned(153, 8)),
	833 => std_logic_vector(to_unsigned(160, 8)),
	834 => std_logic_vector(to_unsigned(165, 8)),
	835 => std_logic_vector(to_unsigned(152, 8)),
	836 => std_logic_vector(to_unsigned(150, 8)),
	837 => std_logic_vector(to_unsigned(155, 8)),
	838 => std_logic_vector(to_unsigned(166, 8)),
	839 => std_logic_vector(to_unsigned(164, 8)),
	840 => std_logic_vector(to_unsigned(165, 8)),
	841 => std_logic_vector(to_unsigned(161, 8)),
	842 => std_logic_vector(to_unsigned(160, 8)),
	843 => std_logic_vector(to_unsigned(166, 8)),
	844 => std_logic_vector(to_unsigned(157, 8)),
	845 => std_logic_vector(to_unsigned(165, 8)),
	846 => std_logic_vector(to_unsigned(160, 8)),
	847 => std_logic_vector(to_unsigned(166, 8)),
	848 => std_logic_vector(to_unsigned(151, 8)),
	849 => std_logic_vector(to_unsigned(163, 8)),
	850 => std_logic_vector(to_unsigned(154, 8)),
	851 => std_logic_vector(to_unsigned(160, 8)),
	852 => std_logic_vector(to_unsigned(160, 8)),
	853 => std_logic_vector(to_unsigned(151, 8)),
	854 => std_logic_vector(to_unsigned(162, 8)),
	855 => std_logic_vector(to_unsigned(166, 8)),
	856 => std_logic_vector(to_unsigned(156, 8)),
	857 => std_logic_vector(to_unsigned(151, 8)),
	858 => std_logic_vector(to_unsigned(152, 8)),
	859 => std_logic_vector(to_unsigned(163, 8)),
	860 => std_logic_vector(to_unsigned(165, 8)),
	861 => std_logic_vector(to_unsigned(161, 8)),
	862 => std_logic_vector(to_unsigned(154, 8)),
	863 => std_logic_vector(to_unsigned(163, 8)),
	864 => std_logic_vector(to_unsigned(154, 8)),
	865 => std_logic_vector(to_unsigned(159, 8)),
	866 => std_logic_vector(to_unsigned(158, 8)),
	867 => std_logic_vector(to_unsigned(154, 8)),
	868 => std_logic_vector(to_unsigned(151, 8)),
	869 => std_logic_vector(to_unsigned(156, 8)),
	870 => std_logic_vector(to_unsigned(164, 8)),
	871 => std_logic_vector(to_unsigned(157, 8)),
	872 => std_logic_vector(to_unsigned(161, 8)),
	873 => std_logic_vector(to_unsigned(162, 8)),
	874 => std_logic_vector(to_unsigned(161, 8)),
	875 => std_logic_vector(to_unsigned(153, 8)),
	876 => std_logic_vector(to_unsigned(165, 8)),
	877 => std_logic_vector(to_unsigned(161, 8)),
	878 => std_logic_vector(to_unsigned(151, 8)),
	879 => std_logic_vector(to_unsigned(156, 8)),
	880 => std_logic_vector(to_unsigned(166, 8)),
	881 => std_logic_vector(to_unsigned(164, 8)),
	882 => std_logic_vector(to_unsigned(158, 8)),
	883 => std_logic_vector(to_unsigned(154, 8)),
	884 => std_logic_vector(to_unsigned(165, 8)),
	885 => std_logic_vector(to_unsigned(161, 8)),
	886 => std_logic_vector(to_unsigned(161, 8)),
	887 => std_logic_vector(to_unsigned(161, 8)),
	888 => std_logic_vector(to_unsigned(162, 8)),
	889 => std_logic_vector(to_unsigned(154, 8)),
	others =>(others =>'0'));

component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_rst         : in  std_logic;
      i_start       : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector (7 downto 0)
      );
end component project_reti_logiche;


begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_rst      	=> tb_rst,
          i_start       => tb_start,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
          o_we 		=> mem_we,
          o_data    	=> mem_i_data
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;


MEM : process(tb_clk)
begin
    if tb_clk'event and tb_clk = '1' then
        if enable_wire = '1' then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
            end if;
        end if;
    end if;
end process;


test : process is
begin
    wait for 55 ns;
    -- wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    -- wait for c_CLOCK_PERIOD;
    -- wait for 100 ns;
    wait for 10 ns;
    tb_rst <= '0';
    -- wait for c_CLOCK_PERIOD;
    -- wait for 100 ns;
    tb_start <= '1';
    -- wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    -- wait for c_CLOCK_PERIOD;
    wait for 10 ns;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;

    assert RAM(890) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(890)))) severity failure;
    assert RAM(891) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(891)))) severity failure;
    assert RAM(892) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(892)))) severity failure;
    assert RAM(893) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(893)))) severity failure;
    assert RAM(894) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(894)))) severity failure;
    assert RAM(895) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(895)))) severity failure;
    assert RAM(896) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(896)))) severity failure;
    assert RAM(897) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(897)))) severity failure;
    assert RAM(898) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(898)))) severity failure;
    assert RAM(899) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(899)))) severity failure;
    assert RAM(900) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(900)))) severity failure;
    assert RAM(901) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(901)))) severity failure;
    assert RAM(902) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(902)))) severity failure;
    assert RAM(903) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(903)))) severity failure;
    assert RAM(904) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(904)))) severity failure;
    assert RAM(905) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(905)))) severity failure;
    assert RAM(906) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(906)))) severity failure;
    assert RAM(907) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(907)))) severity failure;
    assert RAM(908) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(908)))) severity failure;
    assert RAM(909) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(909)))) severity failure;
    assert RAM(910) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(910)))) severity failure;
    assert RAM(911) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(911)))) severity failure;
    assert RAM(912) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(912)))) severity failure;
    assert RAM(913) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(913)))) severity failure;
    assert RAM(914) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(914)))) severity failure;
    assert RAM(915) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(915)))) severity failure;
    assert RAM(916) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(916)))) severity failure;
    assert RAM(917) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(917)))) severity failure;
    assert RAM(918) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(918)))) severity failure;
    assert RAM(919) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(919)))) severity failure;
    assert RAM(920) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(920)))) severity failure;
    assert RAM(921) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(921)))) severity failure;
    assert RAM(922) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(922)))) severity failure;
    assert RAM(923) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(923)))) severity failure;
    assert RAM(924) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(924)))) severity failure;
    assert RAM(925) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(925)))) severity failure;
    assert RAM(926) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(926)))) severity failure;
    assert RAM(927) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(927)))) severity failure;
    assert RAM(928) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(928)))) severity failure;
    assert RAM(929) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(929)))) severity failure;
    assert RAM(930) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(930)))) severity failure;
    assert RAM(931) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(931)))) severity failure;
    assert RAM(932) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(932)))) severity failure;
    assert RAM(933) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(933)))) severity failure;
    assert RAM(934) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(934)))) severity failure;
    assert RAM(935) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(935)))) severity failure;
    assert RAM(936) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(936)))) severity failure;
    assert RAM(937) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(937)))) severity failure;
    assert RAM(938) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(938)))) severity failure;
    assert RAM(939) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(939)))) severity failure;
    assert RAM(940) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(940)))) severity failure;
    assert RAM(941) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(941)))) severity failure;
    assert RAM(942) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(942)))) severity failure;
    assert RAM(943) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(943)))) severity failure;
    assert RAM(944) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(944)))) severity failure;
    assert RAM(945) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(945)))) severity failure;
    assert RAM(946) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(946)))) severity failure;
    assert RAM(947) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(947)))) severity failure;
    assert RAM(948) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(948)))) severity failure;
    assert RAM(949) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(949)))) severity failure;
    assert RAM(950) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(950)))) severity failure;
    assert RAM(951) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(951)))) severity failure;
    assert RAM(952) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(952)))) severity failure;
    assert RAM(953) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(953)))) severity failure;
    assert RAM(954) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(954)))) severity failure;
    assert RAM(955) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(955)))) severity failure;
    assert RAM(956) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(956)))) severity failure;
    assert RAM(957) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(957)))) severity failure;
    assert RAM(958) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(958)))) severity failure;
    assert RAM(959) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(959)))) severity failure;
    assert RAM(960) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(960)))) severity failure;
    assert RAM(961) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(961)))) severity failure;
    assert RAM(962) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(962)))) severity failure;
    assert RAM(963) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(963)))) severity failure;
    assert RAM(964) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(964)))) severity failure;
    assert RAM(965) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(965)))) severity failure;
    assert RAM(966) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(966)))) severity failure;
    assert RAM(967) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(967)))) severity failure;
    assert RAM(968) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(968)))) severity failure;
    assert RAM(969) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(969)))) severity failure;
    assert RAM(970) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(970)))) severity failure;
    assert RAM(971) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(971)))) severity failure;
    assert RAM(972) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(972)))) severity failure;
    assert RAM(973) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(973)))) severity failure;
    assert RAM(974) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(974)))) severity failure;
    assert RAM(975) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(975)))) severity failure;
    assert RAM(976) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(976)))) severity failure;
    assert RAM(977) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(977)))) severity failure;
    assert RAM(978) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(978)))) severity failure;
    assert RAM(979) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(979)))) severity failure;
    assert RAM(980) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(980)))) severity failure;
    assert RAM(981) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(981)))) severity failure;
    assert RAM(982) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(982)))) severity failure;
    assert RAM(983) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(983)))) severity failure;
    assert RAM(984) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(984)))) severity failure;
    assert RAM(985) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(985)))) severity failure;
    assert RAM(986) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(986)))) severity failure;
    assert RAM(987) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(987)))) severity failure;
    assert RAM(988) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(988)))) severity failure;
    assert RAM(989) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(989)))) severity failure;
    assert RAM(990) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(990)))) severity failure;
    assert RAM(991) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(991)))) severity failure;
    assert RAM(992) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(992)))) severity failure;
    assert RAM(993) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(993)))) severity failure;
    assert RAM(994) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(994)))) severity failure;
    assert RAM(995) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(995)))) severity failure;
    assert RAM(996) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(996)))) severity failure;
    assert RAM(997) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(997)))) severity failure;
    assert RAM(998) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(998)))) severity failure;
    assert RAM(999) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(999)))) severity failure;
    assert RAM(1000) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1000)))) severity failure;
    assert RAM(1001) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1001)))) severity failure;
    assert RAM(1002) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1002)))) severity failure;
    assert RAM(1003) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1003)))) severity failure;
    assert RAM(1004) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1004)))) severity failure;
    assert RAM(1005) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1005)))) severity failure;
    assert RAM(1006) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1006)))) severity failure;
    assert RAM(1007) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1007)))) severity failure;
    assert RAM(1008) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1008)))) severity failure;
    assert RAM(1009) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1009)))) severity failure;
    assert RAM(1010) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1010)))) severity failure;
    assert RAM(1011) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1011)))) severity failure;
    assert RAM(1012) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1012)))) severity failure;
    assert RAM(1013) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1013)))) severity failure;
    assert RAM(1014) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1014)))) severity failure;
    assert RAM(1015) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1015)))) severity failure;
    assert RAM(1016) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1016)))) severity failure;
    assert RAM(1017) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1017)))) severity failure;
    assert RAM(1018) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1018)))) severity failure;
    assert RAM(1019) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1019)))) severity failure;
    assert RAM(1020) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1020)))) severity failure;
    assert RAM(1021) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1021)))) severity failure;
    assert RAM(1022) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1022)))) severity failure;
    assert RAM(1023) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1023)))) severity failure;
    assert RAM(1024) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1024)))) severity failure;
    assert RAM(1025) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1025)))) severity failure;
    assert RAM(1026) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1026)))) severity failure;
    assert RAM(1027) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1027)))) severity failure;
    assert RAM(1028) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1028)))) severity failure;
    assert RAM(1029) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1029)))) severity failure;
    assert RAM(1030) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1030)))) severity failure;
    assert RAM(1031) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1031)))) severity failure;
    assert RAM(1032) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1032)))) severity failure;
    assert RAM(1033) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1033)))) severity failure;
    assert RAM(1034) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1034)))) severity failure;
    assert RAM(1035) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1035)))) severity failure;
    assert RAM(1036) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1036)))) severity failure;
    assert RAM(1037) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1037)))) severity failure;
    assert RAM(1038) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1038)))) severity failure;
    assert RAM(1039) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1039)))) severity failure;
    assert RAM(1040) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1040)))) severity failure;
    assert RAM(1041) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1041)))) severity failure;
    assert RAM(1042) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1042)))) severity failure;
    assert RAM(1043) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1043)))) severity failure;
    assert RAM(1044) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1044)))) severity failure;
    assert RAM(1045) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1045)))) severity failure;
    assert RAM(1046) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1046)))) severity failure;
    assert RAM(1047) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1047)))) severity failure;
    assert RAM(1048) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1048)))) severity failure;
    assert RAM(1049) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1049)))) severity failure;
    assert RAM(1050) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1050)))) severity failure;
    assert RAM(1051) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1051)))) severity failure;
    assert RAM(1052) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1052)))) severity failure;
    assert RAM(1053) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1053)))) severity failure;
    assert RAM(1054) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1054)))) severity failure;
    assert RAM(1055) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1055)))) severity failure;
    assert RAM(1056) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1056)))) severity failure;
    assert RAM(1057) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1057)))) severity failure;
    assert RAM(1058) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1058)))) severity failure;
    assert RAM(1059) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1059)))) severity failure;
    assert RAM(1060) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1060)))) severity failure;
    assert RAM(1061) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1061)))) severity failure;
    assert RAM(1062) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1062)))) severity failure;
    assert RAM(1063) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1063)))) severity failure;
    assert RAM(1064) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1064)))) severity failure;
    assert RAM(1065) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1065)))) severity failure;
    assert RAM(1066) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1066)))) severity failure;
    assert RAM(1067) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1067)))) severity failure;
    assert RAM(1068) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1068)))) severity failure;
    assert RAM(1069) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1069)))) severity failure;
    assert RAM(1070) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1070)))) severity failure;
    assert RAM(1071) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1071)))) severity failure;
    assert RAM(1072) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1072)))) severity failure;
    assert RAM(1073) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1073)))) severity failure;
    assert RAM(1074) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1074)))) severity failure;
    assert RAM(1075) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1075)))) severity failure;
    assert RAM(1076) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1076)))) severity failure;
    assert RAM(1077) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1077)))) severity failure;
    assert RAM(1078) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1078)))) severity failure;
    assert RAM(1079) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1079)))) severity failure;
    assert RAM(1080) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1080)))) severity failure;
    assert RAM(1081) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1081)))) severity failure;
    assert RAM(1082) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1082)))) severity failure;
    assert RAM(1083) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1083)))) severity failure;
    assert RAM(1084) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1084)))) severity failure;
    assert RAM(1085) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1085)))) severity failure;
    assert RAM(1086) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1086)))) severity failure;
    assert RAM(1087) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1087)))) severity failure;
    assert RAM(1088) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1088)))) severity failure;
    assert RAM(1089) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1089)))) severity failure;
    assert RAM(1090) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1090)))) severity failure;
    assert RAM(1091) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1091)))) severity failure;
    assert RAM(1092) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1092)))) severity failure;
    assert RAM(1093) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1093)))) severity failure;
    assert RAM(1094) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1094)))) severity failure;
    assert RAM(1095) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1095)))) severity failure;
    assert RAM(1096) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1096)))) severity failure;
    assert RAM(1097) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1097)))) severity failure;
    assert RAM(1098) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1098)))) severity failure;
    assert RAM(1099) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1099)))) severity failure;
    assert RAM(1100) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1100)))) severity failure;
    assert RAM(1101) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1101)))) severity failure;
    assert RAM(1102) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1102)))) severity failure;
    assert RAM(1103) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1103)))) severity failure;
    assert RAM(1104) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1104)))) severity failure;
    assert RAM(1105) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1105)))) severity failure;
    assert RAM(1106) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1106)))) severity failure;
    assert RAM(1107) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1107)))) severity failure;
    assert RAM(1108) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1108)))) severity failure;
    assert RAM(1109) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1109)))) severity failure;
    assert RAM(1110) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1110)))) severity failure;
    assert RAM(1111) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1111)))) severity failure;
    assert RAM(1112) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1112)))) severity failure;
    assert RAM(1113) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1113)))) severity failure;
    assert RAM(1114) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1114)))) severity failure;
    assert RAM(1115) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1115)))) severity failure;
    assert RAM(1116) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1116)))) severity failure;
    assert RAM(1117) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1117)))) severity failure;
    assert RAM(1118) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1118)))) severity failure;
    assert RAM(1119) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1119)))) severity failure;
    assert RAM(1120) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1120)))) severity failure;
    assert RAM(1121) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1121)))) severity failure;
    assert RAM(1122) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1122)))) severity failure;
    assert RAM(1123) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1123)))) severity failure;
    assert RAM(1124) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1124)))) severity failure;
    assert RAM(1125) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1125)))) severity failure;
    assert RAM(1126) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1126)))) severity failure;
    assert RAM(1127) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1127)))) severity failure;
    assert RAM(1128) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1128)))) severity failure;
    assert RAM(1129) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1129)))) severity failure;
    assert RAM(1130) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1130)))) severity failure;
    assert RAM(1131) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1131)))) severity failure;
    assert RAM(1132) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1132)))) severity failure;
    assert RAM(1133) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1133)))) severity failure;
    assert RAM(1134) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1134)))) severity failure;
    assert RAM(1135) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1135)))) severity failure;
    assert RAM(1136) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1136)))) severity failure;
    assert RAM(1137) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1137)))) severity failure;
    assert RAM(1138) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1138)))) severity failure;
    assert RAM(1139) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1139)))) severity failure;
    assert RAM(1140) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1140)))) severity failure;
    assert RAM(1141) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1141)))) severity failure;
    assert RAM(1142) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1142)))) severity failure;
    assert RAM(1143) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1143)))) severity failure;
    assert RAM(1144) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1144)))) severity failure;
    assert RAM(1145) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1145)))) severity failure;
    assert RAM(1146) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1146)))) severity failure;
    assert RAM(1147) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1147)))) severity failure;
    assert RAM(1148) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1148)))) severity failure;
    assert RAM(1149) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1149)))) severity failure;
    assert RAM(1150) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1150)))) severity failure;
    assert RAM(1151) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1151)))) severity failure;
    assert RAM(1152) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1152)))) severity failure;
    assert RAM(1153) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1153)))) severity failure;
    assert RAM(1154) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1154)))) severity failure;
    assert RAM(1155) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1155)))) severity failure;
    assert RAM(1156) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1156)))) severity failure;
    assert RAM(1157) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1157)))) severity failure;
    assert RAM(1158) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1158)))) severity failure;
    assert RAM(1159) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1159)))) severity failure;
    assert RAM(1160) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1160)))) severity failure;
    assert RAM(1161) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1161)))) severity failure;
    assert RAM(1162) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1162)))) severity failure;
    assert RAM(1163) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1163)))) severity failure;
    assert RAM(1164) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1164)))) severity failure;
    assert RAM(1165) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1165)))) severity failure;
    assert RAM(1166) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1166)))) severity failure;
    assert RAM(1167) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1167)))) severity failure;
    assert RAM(1168) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1168)))) severity failure;
    assert RAM(1169) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1169)))) severity failure;
    assert RAM(1170) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1170)))) severity failure;
    assert RAM(1171) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1171)))) severity failure;
    assert RAM(1172) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1172)))) severity failure;
    assert RAM(1173) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1173)))) severity failure;
    assert RAM(1174) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1174)))) severity failure;
    assert RAM(1175) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1175)))) severity failure;
    assert RAM(1176) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1176)))) severity failure;
    assert RAM(1177) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1177)))) severity failure;
    assert RAM(1178) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1178)))) severity failure;
    assert RAM(1179) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1179)))) severity failure;
    assert RAM(1180) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1180)))) severity failure;
    assert RAM(1181) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1181)))) severity failure;
    assert RAM(1182) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1182)))) severity failure;
    assert RAM(1183) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1183)))) severity failure;
    assert RAM(1184) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1184)))) severity failure;
    assert RAM(1185) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1185)))) severity failure;
    assert RAM(1186) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1186)))) severity failure;
    assert RAM(1187) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1187)))) severity failure;
    assert RAM(1188) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1188)))) severity failure;
    assert RAM(1189) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1189)))) severity failure;
    assert RAM(1190) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1190)))) severity failure;
    assert RAM(1191) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1191)))) severity failure;
    assert RAM(1192) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1192)))) severity failure;
    assert RAM(1193) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1193)))) severity failure;
    assert RAM(1194) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1194)))) severity failure;
    assert RAM(1195) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1195)))) severity failure;
    assert RAM(1196) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1196)))) severity failure;
    assert RAM(1197) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1197)))) severity failure;
    assert RAM(1198) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1198)))) severity failure;
    assert RAM(1199) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1199)))) severity failure;
    assert RAM(1200) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1200)))) severity failure;
    assert RAM(1201) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1201)))) severity failure;
    assert RAM(1202) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1202)))) severity failure;
    assert RAM(1203) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1203)))) severity failure;
    assert RAM(1204) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1204)))) severity failure;
    assert RAM(1205) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1205)))) severity failure;
    assert RAM(1206) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1206)))) severity failure;
    assert RAM(1207) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1207)))) severity failure;
    assert RAM(1208) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1208)))) severity failure;
    assert RAM(1209) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1209)))) severity failure;
    assert RAM(1210) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1210)))) severity failure;
    assert RAM(1211) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1211)))) severity failure;
    assert RAM(1212) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1212)))) severity failure;
    assert RAM(1213) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1213)))) severity failure;
    assert RAM(1214) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1214)))) severity failure;
    assert RAM(1215) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1215)))) severity failure;
    assert RAM(1216) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1216)))) severity failure;
    assert RAM(1217) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1217)))) severity failure;
    assert RAM(1218) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1218)))) severity failure;
    assert RAM(1219) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1219)))) severity failure;
    assert RAM(1220) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1220)))) severity failure;
    assert RAM(1221) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1221)))) severity failure;
    assert RAM(1222) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1222)))) severity failure;
    assert RAM(1223) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1223)))) severity failure;
    assert RAM(1224) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1224)))) severity failure;
    assert RAM(1225) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1225)))) severity failure;
    assert RAM(1226) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1226)))) severity failure;
    assert RAM(1227) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1227)))) severity failure;
    assert RAM(1228) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1228)))) severity failure;
    assert RAM(1229) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1229)))) severity failure;
    assert RAM(1230) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1230)))) severity failure;
    assert RAM(1231) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1231)))) severity failure;
    assert RAM(1232) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1232)))) severity failure;
    assert RAM(1233) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1233)))) severity failure;
    assert RAM(1234) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1234)))) severity failure;
    assert RAM(1235) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1235)))) severity failure;
    assert RAM(1236) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1236)))) severity failure;
    assert RAM(1237) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1237)))) severity failure;
    assert RAM(1238) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1238)))) severity failure;
    assert RAM(1239) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1239)))) severity failure;
    assert RAM(1240) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1240)))) severity failure;
    assert RAM(1241) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1241)))) severity failure;
    assert RAM(1242) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1242)))) severity failure;
    assert RAM(1243) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1243)))) severity failure;
    assert RAM(1244) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1244)))) severity failure;
    assert RAM(1245) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1245)))) severity failure;
    assert RAM(1246) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1246)))) severity failure;
    assert RAM(1247) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1247)))) severity failure;
    assert RAM(1248) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1248)))) severity failure;
    assert RAM(1249) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1249)))) severity failure;
    assert RAM(1250) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1250)))) severity failure;
    assert RAM(1251) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1251)))) severity failure;
    assert RAM(1252) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1252)))) severity failure;
    assert RAM(1253) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1253)))) severity failure;
    assert RAM(1254) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1254)))) severity failure;
    assert RAM(1255) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1255)))) severity failure;
    assert RAM(1256) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1256)))) severity failure;
    assert RAM(1257) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1257)))) severity failure;
    assert RAM(1258) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1258)))) severity failure;
    assert RAM(1259) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1259)))) severity failure;
    assert RAM(1260) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1260)))) severity failure;
    assert RAM(1261) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1261)))) severity failure;
    assert RAM(1262) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1262)))) severity failure;
    assert RAM(1263) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1263)))) severity failure;
    assert RAM(1264) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1264)))) severity failure;
    assert RAM(1265) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1265)))) severity failure;
    assert RAM(1266) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1266)))) severity failure;
    assert RAM(1267) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1267)))) severity failure;
    assert RAM(1268) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1268)))) severity failure;
    assert RAM(1269) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1269)))) severity failure;
    assert RAM(1270) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1270)))) severity failure;
    assert RAM(1271) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1271)))) severity failure;
    assert RAM(1272) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1272)))) severity failure;
    assert RAM(1273) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1273)))) severity failure;
    assert RAM(1274) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1274)))) severity failure;
    assert RAM(1275) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1275)))) severity failure;
    assert RAM(1276) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1276)))) severity failure;
    assert RAM(1277) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1277)))) severity failure;
    assert RAM(1278) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1278)))) severity failure;
    assert RAM(1279) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1279)))) severity failure;
    assert RAM(1280) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1280)))) severity failure;
    assert RAM(1281) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1281)))) severity failure;
    assert RAM(1282) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1282)))) severity failure;
    assert RAM(1283) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1283)))) severity failure;
    assert RAM(1284) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1284)))) severity failure;
    assert RAM(1285) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1285)))) severity failure;
    assert RAM(1286) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1286)))) severity failure;
    assert RAM(1287) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1287)))) severity failure;
    assert RAM(1288) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1288)))) severity failure;
    assert RAM(1289) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1289)))) severity failure;
    assert RAM(1290) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1290)))) severity failure;
    assert RAM(1291) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1291)))) severity failure;
    assert RAM(1292) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1292)))) severity failure;
    assert RAM(1293) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1293)))) severity failure;
    assert RAM(1294) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1294)))) severity failure;
    assert RAM(1295) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1295)))) severity failure;
    assert RAM(1296) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1296)))) severity failure;
    assert RAM(1297) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1297)))) severity failure;
    assert RAM(1298) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1298)))) severity failure;
    assert RAM(1299) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1299)))) severity failure;
    assert RAM(1300) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1300)))) severity failure;
    assert RAM(1301) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1301)))) severity failure;
    assert RAM(1302) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1302)))) severity failure;
    assert RAM(1303) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1303)))) severity failure;
    assert RAM(1304) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1304)))) severity failure;
    assert RAM(1305) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1305)))) severity failure;
    assert RAM(1306) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1306)))) severity failure;
    assert RAM(1307) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1307)))) severity failure;
    assert RAM(1308) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1308)))) severity failure;
    assert RAM(1309) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1309)))) severity failure;
    assert RAM(1310) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1310)))) severity failure;
    assert RAM(1311) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1311)))) severity failure;
    assert RAM(1312) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1312)))) severity failure;
    assert RAM(1313) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1313)))) severity failure;
    assert RAM(1314) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1314)))) severity failure;
    assert RAM(1315) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1315)))) severity failure;
    assert RAM(1316) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1316)))) severity failure;
    assert RAM(1317) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1317)))) severity failure;
    assert RAM(1318) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1318)))) severity failure;
    assert RAM(1319) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1319)))) severity failure;
    assert RAM(1320) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1320)))) severity failure;
    assert RAM(1321) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1321)))) severity failure;
    assert RAM(1322) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1322)))) severity failure;
    assert RAM(1323) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1323)))) severity failure;
    assert RAM(1324) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1324)))) severity failure;
    assert RAM(1325) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1325)))) severity failure;
    assert RAM(1326) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1326)))) severity failure;
    assert RAM(1327) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1327)))) severity failure;
    assert RAM(1328) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1328)))) severity failure;
    assert RAM(1329) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1329)))) severity failure;
    assert RAM(1330) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1330)))) severity failure;
    assert RAM(1331) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1331)))) severity failure;
    assert RAM(1332) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1332)))) severity failure;
    assert RAM(1333) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1333)))) severity failure;
    assert RAM(1334) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1334)))) severity failure;
    assert RAM(1335) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1335)))) severity failure;
    assert RAM(1336) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1336)))) severity failure;
    assert RAM(1337) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1337)))) severity failure;
    assert RAM(1338) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1338)))) severity failure;
    assert RAM(1339) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1339)))) severity failure;
    assert RAM(1340) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1340)))) severity failure;
    assert RAM(1341) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1341)))) severity failure;
    assert RAM(1342) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1342)))) severity failure;
    assert RAM(1343) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1343)))) severity failure;
    assert RAM(1344) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1344)))) severity failure;
    assert RAM(1345) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1345)))) severity failure;
    assert RAM(1346) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1346)))) severity failure;
    assert RAM(1347) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1347)))) severity failure;
    assert RAM(1348) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1348)))) severity failure;
    assert RAM(1349) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1349)))) severity failure;
    assert RAM(1350) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1350)))) severity failure;
    assert RAM(1351) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1351)))) severity failure;
    assert RAM(1352) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1352)))) severity failure;
    assert RAM(1353) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1353)))) severity failure;
    assert RAM(1354) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1354)))) severity failure;
    assert RAM(1355) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1355)))) severity failure;
    assert RAM(1356) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1356)))) severity failure;
    assert RAM(1357) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1357)))) severity failure;
    assert RAM(1358) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1358)))) severity failure;
    assert RAM(1359) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1359)))) severity failure;
    assert RAM(1360) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1360)))) severity failure;
    assert RAM(1361) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1361)))) severity failure;
    assert RAM(1362) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1362)))) severity failure;
    assert RAM(1363) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1363)))) severity failure;
    assert RAM(1364) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1364)))) severity failure;
    assert RAM(1365) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1365)))) severity failure;
    assert RAM(1366) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1366)))) severity failure;
    assert RAM(1367) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1367)))) severity failure;
    assert RAM(1368) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1368)))) severity failure;
    assert RAM(1369) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1369)))) severity failure;
    assert RAM(1370) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1370)))) severity failure;
    assert RAM(1371) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1371)))) severity failure;
    assert RAM(1372) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1372)))) severity failure;
    assert RAM(1373) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1373)))) severity failure;
    assert RAM(1374) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1374)))) severity failure;
    assert RAM(1375) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1375)))) severity failure;
    assert RAM(1376) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1376)))) severity failure;
    assert RAM(1377) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1377)))) severity failure;
    assert RAM(1378) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1378)))) severity failure;
    assert RAM(1379) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1379)))) severity failure;
    assert RAM(1380) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1380)))) severity failure;
    assert RAM(1381) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1381)))) severity failure;
    assert RAM(1382) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1382)))) severity failure;
    assert RAM(1383) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1383)))) severity failure;
    assert RAM(1384) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1384)))) severity failure;
    assert RAM(1385) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1385)))) severity failure;
    assert RAM(1386) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1386)))) severity failure;
    assert RAM(1387) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1387)))) severity failure;
    assert RAM(1388) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1388)))) severity failure;
    assert RAM(1389) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1389)))) severity failure;
    assert RAM(1390) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1390)))) severity failure;
    assert RAM(1391) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1391)))) severity failure;
    assert RAM(1392) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1392)))) severity failure;
    assert RAM(1393) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1393)))) severity failure;
    assert RAM(1394) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1394)))) severity failure;
    assert RAM(1395) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1395)))) severity failure;
    assert RAM(1396) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1396)))) severity failure;
    assert RAM(1397) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1397)))) severity failure;
    assert RAM(1398) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1398)))) severity failure;
    assert RAM(1399) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1399)))) severity failure;
    assert RAM(1400) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1400)))) severity failure;
    assert RAM(1401) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1401)))) severity failure;
    assert RAM(1402) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1402)))) severity failure;
    assert RAM(1403) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1403)))) severity failure;
    assert RAM(1404) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1404)))) severity failure;
    assert RAM(1405) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1405)))) severity failure;
    assert RAM(1406) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1406)))) severity failure;
    assert RAM(1407) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1407)))) severity failure;
    assert RAM(1408) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1408)))) severity failure;
    assert RAM(1409) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1409)))) severity failure;
    assert RAM(1410) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1410)))) severity failure;
    assert RAM(1411) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1411)))) severity failure;
    assert RAM(1412) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1412)))) severity failure;
    assert RAM(1413) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1413)))) severity failure;
    assert RAM(1414) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1414)))) severity failure;
    assert RAM(1415) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1415)))) severity failure;
    assert RAM(1416) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1416)))) severity failure;
    assert RAM(1417) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1417)))) severity failure;
    assert RAM(1418) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1418)))) severity failure;
    assert RAM(1419) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1419)))) severity failure;
    assert RAM(1420) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1420)))) severity failure;
    assert RAM(1421) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1421)))) severity failure;
    assert RAM(1422) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1422)))) severity failure;
    assert RAM(1423) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1423)))) severity failure;
    assert RAM(1424) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1424)))) severity failure;
    assert RAM(1425) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1425)))) severity failure;
    assert RAM(1426) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1426)))) severity failure;
    assert RAM(1427) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1427)))) severity failure;
    assert RAM(1428) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1428)))) severity failure;
    assert RAM(1429) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1429)))) severity failure;
    assert RAM(1430) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1430)))) severity failure;
    assert RAM(1431) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1431)))) severity failure;
    assert RAM(1432) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1432)))) severity failure;
    assert RAM(1433) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1433)))) severity failure;
    assert RAM(1434) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1434)))) severity failure;
    assert RAM(1435) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1435)))) severity failure;
    assert RAM(1436) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1436)))) severity failure;
    assert RAM(1437) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1437)))) severity failure;
    assert RAM(1438) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1438)))) severity failure;
    assert RAM(1439) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1439)))) severity failure;
    assert RAM(1440) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1440)))) severity failure;
    assert RAM(1441) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1441)))) severity failure;
    assert RAM(1442) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1442)))) severity failure;
    assert RAM(1443) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1443)))) severity failure;
    assert RAM(1444) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1444)))) severity failure;
    assert RAM(1445) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1445)))) severity failure;
    assert RAM(1446) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1446)))) severity failure;
    assert RAM(1447) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1447)))) severity failure;
    assert RAM(1448) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1448)))) severity failure;
    assert RAM(1449) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1449)))) severity failure;
    assert RAM(1450) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1450)))) severity failure;
    assert RAM(1451) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1451)))) severity failure;
    assert RAM(1452) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1452)))) severity failure;
    assert RAM(1453) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1453)))) severity failure;
    assert RAM(1454) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1454)))) severity failure;
    assert RAM(1455) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1455)))) severity failure;
    assert RAM(1456) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1456)))) severity failure;
    assert RAM(1457) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1457)))) severity failure;
    assert RAM(1458) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1458)))) severity failure;
    assert RAM(1459) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1459)))) severity failure;
    assert RAM(1460) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1460)))) severity failure;
    assert RAM(1461) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1461)))) severity failure;
    assert RAM(1462) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1462)))) severity failure;
    assert RAM(1463) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1463)))) severity failure;
    assert RAM(1464) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1464)))) severity failure;
    assert RAM(1465) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1465)))) severity failure;
    assert RAM(1466) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1466)))) severity failure;
    assert RAM(1467) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1467)))) severity failure;
    assert RAM(1468) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1468)))) severity failure;
    assert RAM(1469) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1469)))) severity failure;
    assert RAM(1470) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1470)))) severity failure;
    assert RAM(1471) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1471)))) severity failure;
    assert RAM(1472) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1472)))) severity failure;
    assert RAM(1473) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1473)))) severity failure;
    assert RAM(1474) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1474)))) severity failure;
    assert RAM(1475) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1475)))) severity failure;
    assert RAM(1476) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1476)))) severity failure;
    assert RAM(1477) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1477)))) severity failure;
    assert RAM(1478) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1478)))) severity failure;
    assert RAM(1479) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1479)))) severity failure;
    assert RAM(1480) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1480)))) severity failure;
    assert RAM(1481) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1481)))) severity failure;
    assert RAM(1482) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1482)))) severity failure;
    assert RAM(1483) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1483)))) severity failure;
    assert RAM(1484) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1484)))) severity failure;
    assert RAM(1485) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1485)))) severity failure;
    assert RAM(1486) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1486)))) severity failure;
    assert RAM(1487) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1487)))) severity failure;
    assert RAM(1488) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1488)))) severity failure;
    assert RAM(1489) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1489)))) severity failure;
    assert RAM(1490) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1490)))) severity failure;
    assert RAM(1491) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1491)))) severity failure;
    assert RAM(1492) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1492)))) severity failure;
    assert RAM(1493) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1493)))) severity failure;
    assert RAM(1494) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1494)))) severity failure;
    assert RAM(1495) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1495)))) severity failure;
    assert RAM(1496) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1496)))) severity failure;
    assert RAM(1497) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1497)))) severity failure;
    assert RAM(1498) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1498)))) severity failure;
    assert RAM(1499) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1499)))) severity failure;
    assert RAM(1500) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1500)))) severity failure;
    assert RAM(1501) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1501)))) severity failure;
    assert RAM(1502) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1502)))) severity failure;
    assert RAM(1503) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1503)))) severity failure;
    assert RAM(1504) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1504)))) severity failure;
    assert RAM(1505) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1505)))) severity failure;
    assert RAM(1506) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1506)))) severity failure;
    assert RAM(1507) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1507)))) severity failure;
    assert RAM(1508) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1508)))) severity failure;
    assert RAM(1509) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1509)))) severity failure;
    assert RAM(1510) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1510)))) severity failure;
    assert RAM(1511) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1511)))) severity failure;
    assert RAM(1512) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1512)))) severity failure;
    assert RAM(1513) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1513)))) severity failure;
    assert RAM(1514) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1514)))) severity failure;
    assert RAM(1515) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1515)))) severity failure;
    assert RAM(1516) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1516)))) severity failure;
    assert RAM(1517) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1517)))) severity failure;
    assert RAM(1518) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1518)))) severity failure;
    assert RAM(1519) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1519)))) severity failure;
    assert RAM(1520) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1520)))) severity failure;
    assert RAM(1521) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1521)))) severity failure;
    assert RAM(1522) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1522)))) severity failure;
    assert RAM(1523) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1523)))) severity failure;
    assert RAM(1524) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1524)))) severity failure;
    assert RAM(1525) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1525)))) severity failure;
    assert RAM(1526) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1526)))) severity failure;
    assert RAM(1527) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1527)))) severity failure;
    assert RAM(1528) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1528)))) severity failure;
    assert RAM(1529) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1529)))) severity failure;
    assert RAM(1530) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1530)))) severity failure;
    assert RAM(1531) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1531)))) severity failure;
    assert RAM(1532) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1532)))) severity failure;
    assert RAM(1533) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1533)))) severity failure;
    assert RAM(1534) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1534)))) severity failure;
    assert RAM(1535) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1535)))) severity failure;
    assert RAM(1536) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1536)))) severity failure;
    assert RAM(1537) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1537)))) severity failure;
    assert RAM(1538) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1538)))) severity failure;
    assert RAM(1539) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1539)))) severity failure;
    assert RAM(1540) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1540)))) severity failure;
    assert RAM(1541) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1541)))) severity failure;
    assert RAM(1542) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1542)))) severity failure;
    assert RAM(1543) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1543)))) severity failure;
    assert RAM(1544) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1544)))) severity failure;
    assert RAM(1545) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1545)))) severity failure;
    assert RAM(1546) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1546)))) severity failure;
    assert RAM(1547) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1547)))) severity failure;
    assert RAM(1548) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1548)))) severity failure;
    assert RAM(1549) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1549)))) severity failure;
    assert RAM(1550) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1550)))) severity failure;
    assert RAM(1551) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1551)))) severity failure;
    assert RAM(1552) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1552)))) severity failure;
    assert RAM(1553) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1553)))) severity failure;
    assert RAM(1554) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1554)))) severity failure;
    assert RAM(1555) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1555)))) severity failure;
    assert RAM(1556) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1556)))) severity failure;
    assert RAM(1557) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1557)))) severity failure;
    assert RAM(1558) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1558)))) severity failure;
    assert RAM(1559) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1559)))) severity failure;
    assert RAM(1560) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1560)))) severity failure;
    assert RAM(1561) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1561)))) severity failure;
    assert RAM(1562) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1562)))) severity failure;
    assert RAM(1563) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1563)))) severity failure;
    assert RAM(1564) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1564)))) severity failure;
    assert RAM(1565) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1565)))) severity failure;
    assert RAM(1566) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1566)))) severity failure;
    assert RAM(1567) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1567)))) severity failure;
    assert RAM(1568) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1568)))) severity failure;
    assert RAM(1569) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1569)))) severity failure;
    assert RAM(1570) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1570)))) severity failure;
    assert RAM(1571) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1571)))) severity failure;
    assert RAM(1572) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1572)))) severity failure;
    assert RAM(1573) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1573)))) severity failure;
    assert RAM(1574) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1574)))) severity failure;
    assert RAM(1575) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1575)))) severity failure;
    assert RAM(1576) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1576)))) severity failure;
    assert RAM(1577) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1577)))) severity failure;
    assert RAM(1578) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1578)))) severity failure;
    assert RAM(1579) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1579)))) severity failure;
    assert RAM(1580) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1580)))) severity failure;
    assert RAM(1581) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1581)))) severity failure;
    assert RAM(1582) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1582)))) severity failure;
    assert RAM(1583) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1583)))) severity failure;
    assert RAM(1584) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1584)))) severity failure;
    assert RAM(1585) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1585)))) severity failure;
    assert RAM(1586) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1586)))) severity failure;
    assert RAM(1587) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1587)))) severity failure;
    assert RAM(1588) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1588)))) severity failure;
    assert RAM(1589) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1589)))) severity failure;
    assert RAM(1590) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1590)))) severity failure;
    assert RAM(1591) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1591)))) severity failure;
    assert RAM(1592) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1592)))) severity failure;
    assert RAM(1593) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1593)))) severity failure;
    assert RAM(1594) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1594)))) severity failure;
    assert RAM(1595) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1595)))) severity failure;
    assert RAM(1596) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1596)))) severity failure;
    assert RAM(1597) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1597)))) severity failure;
    assert RAM(1598) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1598)))) severity failure;
    assert RAM(1599) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1599)))) severity failure;
    assert RAM(1600) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1600)))) severity failure;
    assert RAM(1601) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1601)))) severity failure;
    assert RAM(1602) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1602)))) severity failure;
    assert RAM(1603) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1603)))) severity failure;
    assert RAM(1604) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1604)))) severity failure;
    assert RAM(1605) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1605)))) severity failure;
    assert RAM(1606) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1606)))) severity failure;
    assert RAM(1607) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1607)))) severity failure;
    assert RAM(1608) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1608)))) severity failure;
    assert RAM(1609) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1609)))) severity failure;
    assert RAM(1610) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1610)))) severity failure;
    assert RAM(1611) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1611)))) severity failure;
    assert RAM(1612) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1612)))) severity failure;
    assert RAM(1613) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1613)))) severity failure;
    assert RAM(1614) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1614)))) severity failure;
    assert RAM(1615) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1615)))) severity failure;
    assert RAM(1616) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1616)))) severity failure;
    assert RAM(1617) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1617)))) severity failure;
    assert RAM(1618) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1618)))) severity failure;
    assert RAM(1619) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1619)))) severity failure;
    assert RAM(1620) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1620)))) severity failure;
    assert RAM(1621) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1621)))) severity failure;
    assert RAM(1622) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1622)))) severity failure;
    assert RAM(1623) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1623)))) severity failure;
    assert RAM(1624) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1624)))) severity failure;
    assert RAM(1625) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1625)))) severity failure;
    assert RAM(1626) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1626)))) severity failure;
    assert RAM(1627) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1627)))) severity failure;
    assert RAM(1628) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1628)))) severity failure;
    assert RAM(1629) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1629)))) severity failure;
    assert RAM(1630) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1630)))) severity failure;
    assert RAM(1631) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1631)))) severity failure;
    assert RAM(1632) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1632)))) severity failure;
    assert RAM(1633) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1633)))) severity failure;
    assert RAM(1634) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1634)))) severity failure;
    assert RAM(1635) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1635)))) severity failure;
    assert RAM(1636) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1636)))) severity failure;
    assert RAM(1637) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1637)))) severity failure;
    assert RAM(1638) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1638)))) severity failure;
    assert RAM(1639) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1639)))) severity failure;
    assert RAM(1640) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1640)))) severity failure;
    assert RAM(1641) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1641)))) severity failure;
    assert RAM(1642) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1642)))) severity failure;
    assert RAM(1643) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1643)))) severity failure;
    assert RAM(1644) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1644)))) severity failure;
    assert RAM(1645) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1645)))) severity failure;
    assert RAM(1646) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1646)))) severity failure;
    assert RAM(1647) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1647)))) severity failure;
    assert RAM(1648) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1648)))) severity failure;
    assert RAM(1649) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1649)))) severity failure;
    assert RAM(1650) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1650)))) severity failure;
    assert RAM(1651) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1651)))) severity failure;
    assert RAM(1652) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1652)))) severity failure;
    assert RAM(1653) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1653)))) severity failure;
    assert RAM(1654) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1654)))) severity failure;
    assert RAM(1655) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1655)))) severity failure;
    assert RAM(1656) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1656)))) severity failure;
    assert RAM(1657) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1657)))) severity failure;
    assert RAM(1658) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1658)))) severity failure;
    assert RAM(1659) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1659)))) severity failure;
    assert RAM(1660) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1660)))) severity failure;
    assert RAM(1661) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1661)))) severity failure;
    assert RAM(1662) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1662)))) severity failure;
    assert RAM(1663) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1663)))) severity failure;
    assert RAM(1664) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1664)))) severity failure;
    assert RAM(1665) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1665)))) severity failure;
    assert RAM(1666) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1666)))) severity failure;
    assert RAM(1667) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1667)))) severity failure;
    assert RAM(1668) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1668)))) severity failure;
    assert RAM(1669) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1669)))) severity failure;
    assert RAM(1670) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1670)))) severity failure;
    assert RAM(1671) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1671)))) severity failure;
    assert RAM(1672) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1672)))) severity failure;
    assert RAM(1673) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1673)))) severity failure;
    assert RAM(1674) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1674)))) severity failure;
    assert RAM(1675) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1675)))) severity failure;
    assert RAM(1676) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1676)))) severity failure;
    assert RAM(1677) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1677)))) severity failure;
    assert RAM(1678) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1678)))) severity failure;
    assert RAM(1679) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1679)))) severity failure;
    assert RAM(1680) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1680)))) severity failure;
    assert RAM(1681) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1681)))) severity failure;
    assert RAM(1682) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1682)))) severity failure;
    assert RAM(1683) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1683)))) severity failure;
    assert RAM(1684) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1684)))) severity failure;
    assert RAM(1685) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1685)))) severity failure;
    assert RAM(1686) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1686)))) severity failure;
    assert RAM(1687) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1687)))) severity failure;
    assert RAM(1688) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1688)))) severity failure;
    assert RAM(1689) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1689)))) severity failure;
    assert RAM(1690) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1690)))) severity failure;
    assert RAM(1691) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1691)))) severity failure;
    assert RAM(1692) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1692)))) severity failure;
    assert RAM(1693) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1693)))) severity failure;
    assert RAM(1694) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1694)))) severity failure;
    assert RAM(1695) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1695)))) severity failure;
    assert RAM(1696) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1696)))) severity failure;
    assert RAM(1697) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1697)))) severity failure;
    assert RAM(1698) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1698)))) severity failure;
    assert RAM(1699) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1699)))) severity failure;
    assert RAM(1700) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1700)))) severity failure;
    assert RAM(1701) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1701)))) severity failure;
    assert RAM(1702) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1702)))) severity failure;
    assert RAM(1703) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1703)))) severity failure;
    assert RAM(1704) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1704)))) severity failure;
    assert RAM(1705) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1705)))) severity failure;
    assert RAM(1706) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1706)))) severity failure;
    assert RAM(1707) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1707)))) severity failure;
    assert RAM(1708) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1708)))) severity failure;
    assert RAM(1709) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1709)))) severity failure;
    assert RAM(1710) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1710)))) severity failure;
    assert RAM(1711) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1711)))) severity failure;
    assert RAM(1712) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1712)))) severity failure;
    assert RAM(1713) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1713)))) severity failure;
    assert RAM(1714) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(1714)))) severity failure;
    assert RAM(1715) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1715)))) severity failure;
    assert RAM(1716) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1716)))) severity failure;
    assert RAM(1717) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1717)))) severity failure;
    assert RAM(1718) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1718)))) severity failure;
    assert RAM(1719) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1719)))) severity failure;
    assert RAM(1720) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1720)))) severity failure;
    assert RAM(1721) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1721)))) severity failure;
    assert RAM(1722) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1722)))) severity failure;
    assert RAM(1723) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1723)))) severity failure;
    assert RAM(1724) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected 16 found " & integer'image(to_integer(unsigned(RAM(1724)))) severity failure;
    assert RAM(1725) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(1725)))) severity failure;
    assert RAM(1726) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1726)))) severity failure;
    assert RAM(1727) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1727)))) severity failure;
    assert RAM(1728) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1728)))) severity failure;
    assert RAM(1729) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1729)))) severity failure;
    assert RAM(1730) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1730)))) severity failure;
    assert RAM(1731) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1731)))) severity failure;
    assert RAM(1732) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1732)))) severity failure;
    assert RAM(1733) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1733)))) severity failure;
    assert RAM(1734) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1734)))) severity failure;
    assert RAM(1735) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1735)))) severity failure;
    assert RAM(1736) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1736)))) severity failure;
    assert RAM(1737) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1737)))) severity failure;
    assert RAM(1738) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1738)))) severity failure;
    assert RAM(1739) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1739)))) severity failure;
    assert RAM(1740) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(1740)))) severity failure;
    assert RAM(1741) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1741)))) severity failure;
    assert RAM(1742) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1742)))) severity failure;
    assert RAM(1743) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1743)))) severity failure;
    assert RAM(1744) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1744)))) severity failure;
    assert RAM(1745) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1745)))) severity failure;
    assert RAM(1746) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected 48 found " & integer'image(to_integer(unsigned(RAM(1746)))) severity failure;
    assert RAM(1747) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1747)))) severity failure;
    assert RAM(1748) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1748)))) severity failure;
    assert RAM(1749) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1749)))) severity failure;
    assert RAM(1750) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1750)))) severity failure;
    assert RAM(1751) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(1751)))) severity failure;
    assert RAM(1752) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1752)))) severity failure;
    assert RAM(1753) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(1753)))) severity failure;
    assert RAM(1754) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1754)))) severity failure;
    assert RAM(1755) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1755)))) severity failure;
    assert RAM(1756) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1756)))) severity failure;
    assert RAM(1757) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1757)))) severity failure;
    assert RAM(1758) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1758)))) severity failure;
    assert RAM(1759) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(1759)))) severity failure;
    assert RAM(1760) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1760)))) severity failure;
    assert RAM(1761) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1761)))) severity failure;
    assert RAM(1762) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1762)))) severity failure;
    assert RAM(1763) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(1763)))) severity failure;
    assert RAM(1764) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1764)))) severity failure;
    assert RAM(1765) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1765)))) severity failure;
    assert RAM(1766) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(1766)))) severity failure;
    assert RAM(1767) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(1767)))) severity failure;
    assert RAM(1768) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1768)))) severity failure;
    assert RAM(1769) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected 240 found " & integer'image(to_integer(unsigned(RAM(1769)))) severity failure;
    assert RAM(1770) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected 144 found " & integer'image(to_integer(unsigned(RAM(1770)))) severity failure;
    assert RAM(1771) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1771)))) severity failure;
    assert RAM(1772) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(1772)))) severity failure;
    assert RAM(1773) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1773)))) severity failure;
    assert RAM(1774) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1774)))) severity failure;
    assert RAM(1775) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(1775)))) severity failure;
    assert RAM(1776) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected 208 found " & integer'image(to_integer(unsigned(RAM(1776)))) severity failure;
    assert RAM(1777) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected 80 found " & integer'image(to_integer(unsigned(RAM(1777)))) severity failure;

    assert false report "Simulation Ended! TEST PASSATO" severity failure;
end process test;

end shlev4tb;
