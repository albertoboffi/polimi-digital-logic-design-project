-------------------------------------------------------------------------------
--
-- Final examination - Digital Logic Design
-- Alberto Boffi - Politecnico di Milano, AY 2020/21
-- TEST MODULE: Consecutive images
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity consimg_tb is
end consimg_tb;

architecture consimgtb of consimg_tb is
constant c_CLOCK_PERIOD         : time := 15 ns;
signal   tb_done                : std_logic;
signal   mem_address            : std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst                 : std_logic := '0';
signal   tb_start               : std_logic := '0';
signal   tb_clk                 : std_logic := '0';
signal   mem_o_data,mem_i_data  : std_logic_vector (7 downto 0);
signal   enable_wire            : std_logic;
signal   mem_we                 : std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);

signal RAM: ram_type :=
	(0 => std_logic_vector(to_unsigned(127, 8)),
	1 => std_logic_vector(to_unsigned(3, 8)),
	2 => std_logic_vector(to_unsigned(108, 8)),
	3 => std_logic_vector(to_unsigned(109, 8)),
	4 => std_logic_vector(to_unsigned(109, 8)),
	5 => std_logic_vector(to_unsigned(106, 8)),
	6 => std_logic_vector(to_unsigned(102, 8)),
	7 => std_logic_vector(to_unsigned(110, 8)),
	8 => std_logic_vector(to_unsigned(103, 8)),
	9 => std_logic_vector(to_unsigned(108, 8)),
	10 => std_logic_vector(to_unsigned(101, 8)),
	11 => std_logic_vector(to_unsigned(107, 8)),
	12 => std_logic_vector(to_unsigned(99, 8)),
	13 => std_logic_vector(to_unsigned(108, 8)),
	14 => std_logic_vector(to_unsigned(109, 8)),
	15 => std_logic_vector(to_unsigned(112, 8)),
	16 => std_logic_vector(to_unsigned(100, 8)),
	17 => std_logic_vector(to_unsigned(100, 8)),
	18 => std_logic_vector(to_unsigned(101, 8)),
	19 => std_logic_vector(to_unsigned(99, 8)),
	20 => std_logic_vector(to_unsigned(100, 8)),
	21 => std_logic_vector(to_unsigned(111, 8)),
	22 => std_logic_vector(to_unsigned(106, 8)),
	23 => std_logic_vector(to_unsigned(102, 8)),
	24 => std_logic_vector(to_unsigned(99, 8)),
	25 => std_logic_vector(to_unsigned(105, 8)),
	26 => std_logic_vector(to_unsigned(105, 8)),
	27 => std_logic_vector(to_unsigned(110, 8)),
	28 => std_logic_vector(to_unsigned(109, 8)),
	29 => std_logic_vector(to_unsigned(109, 8)),
	30 => std_logic_vector(to_unsigned(106, 8)),
	31 => std_logic_vector(to_unsigned(107, 8)),
	32 => std_logic_vector(to_unsigned(101, 8)),
	33 => std_logic_vector(to_unsigned(103, 8)),
	34 => std_logic_vector(to_unsigned(104, 8)),
	35 => std_logic_vector(to_unsigned(104, 8)),
	36 => std_logic_vector(to_unsigned(103, 8)),
	37 => std_logic_vector(to_unsigned(104, 8)),
	38 => std_logic_vector(to_unsigned(102, 8)),
	39 => std_logic_vector(to_unsigned(103, 8)),
	40 => std_logic_vector(to_unsigned(104, 8)),
	41 => std_logic_vector(to_unsigned(106, 8)),
	42 => std_logic_vector(to_unsigned(112, 8)),
	43 => std_logic_vector(to_unsigned(107, 8)),
	44 => std_logic_vector(to_unsigned(99, 8)),
	45 => std_logic_vector(to_unsigned(107, 8)),
	46 => std_logic_vector(to_unsigned(99, 8)),
	47 => std_logic_vector(to_unsigned(112, 8)),
	48 => std_logic_vector(to_unsigned(107, 8)),
	49 => std_logic_vector(to_unsigned(110, 8)),
	50 => std_logic_vector(to_unsigned(104, 8)),
	51 => std_logic_vector(to_unsigned(104, 8)),
	52 => std_logic_vector(to_unsigned(112, 8)),
	53 => std_logic_vector(to_unsigned(112, 8)),
	54 => std_logic_vector(to_unsigned(109, 8)),
	55 => std_logic_vector(to_unsigned(111, 8)),
	56 => std_logic_vector(to_unsigned(105, 8)),
	57 => std_logic_vector(to_unsigned(107, 8)),
	58 => std_logic_vector(to_unsigned(106, 8)),
	59 => std_logic_vector(to_unsigned(101, 8)),
	60 => std_logic_vector(to_unsigned(106, 8)),
	61 => std_logic_vector(to_unsigned(105, 8)),
	62 => std_logic_vector(to_unsigned(101, 8)),
	63 => std_logic_vector(to_unsigned(105, 8)),
	64 => std_logic_vector(to_unsigned(101, 8)),
	65 => std_logic_vector(to_unsigned(104, 8)),
	66 => std_logic_vector(to_unsigned(105, 8)),
	67 => std_logic_vector(to_unsigned(111, 8)),
	68 => std_logic_vector(to_unsigned(111, 8)),
	69 => std_logic_vector(to_unsigned(108, 8)),
	70 => std_logic_vector(to_unsigned(101, 8)),
	71 => std_logic_vector(to_unsigned(101, 8)),
	72 => std_logic_vector(to_unsigned(99, 8)),
	73 => std_logic_vector(to_unsigned(104, 8)),
	74 => std_logic_vector(to_unsigned(110, 8)),
	75 => std_logic_vector(to_unsigned(111, 8)),
	76 => std_logic_vector(to_unsigned(104, 8)),
	77 => std_logic_vector(to_unsigned(99, 8)),
	78 => std_logic_vector(to_unsigned(109, 8)),
	79 => std_logic_vector(to_unsigned(111, 8)),
	80 => std_logic_vector(to_unsigned(99, 8)),
	81 => std_logic_vector(to_unsigned(102, 8)),
	82 => std_logic_vector(to_unsigned(104, 8)),
	83 => std_logic_vector(to_unsigned(107, 8)),
	84 => std_logic_vector(to_unsigned(103, 8)),
	85 => std_logic_vector(to_unsigned(109, 8)),
	86 => std_logic_vector(to_unsigned(112, 8)),
	87 => std_logic_vector(to_unsigned(111, 8)),
	88 => std_logic_vector(to_unsigned(107, 8)),
	89 => std_logic_vector(to_unsigned(106, 8)),
	90 => std_logic_vector(to_unsigned(107, 8)),
	91 => std_logic_vector(to_unsigned(112, 8)),
	92 => std_logic_vector(to_unsigned(99, 8)),
	93 => std_logic_vector(to_unsigned(99, 8)),
	94 => std_logic_vector(to_unsigned(110, 8)),
	95 => std_logic_vector(to_unsigned(104, 8)),
	96 => std_logic_vector(to_unsigned(110, 8)),
	97 => std_logic_vector(to_unsigned(109, 8)),
	98 => std_logic_vector(to_unsigned(101, 8)),
	99 => std_logic_vector(to_unsigned(104, 8)),
	100 => std_logic_vector(to_unsigned(105, 8)),
	101 => std_logic_vector(to_unsigned(111, 8)),
	102 => std_logic_vector(to_unsigned(107, 8)),
	103 => std_logic_vector(to_unsigned(111, 8)),
	104 => std_logic_vector(to_unsigned(111, 8)),
	105 => std_logic_vector(to_unsigned(99, 8)),
	106 => std_logic_vector(to_unsigned(111, 8)),
	107 => std_logic_vector(to_unsigned(105, 8)),
	108 => std_logic_vector(to_unsigned(99, 8)),
	109 => std_logic_vector(to_unsigned(105, 8)),
	110 => std_logic_vector(to_unsigned(100, 8)),
	111 => std_logic_vector(to_unsigned(111, 8)),
	112 => std_logic_vector(to_unsigned(99, 8)),
	113 => std_logic_vector(to_unsigned(104, 8)),
	114 => std_logic_vector(to_unsigned(106, 8)),
	115 => std_logic_vector(to_unsigned(100, 8)),
	116 => std_logic_vector(to_unsigned(103, 8)),
	117 => std_logic_vector(to_unsigned(103, 8)),
	118 => std_logic_vector(to_unsigned(109, 8)),
	119 => std_logic_vector(to_unsigned(99, 8)),
	120 => std_logic_vector(to_unsigned(101, 8)),
	121 => std_logic_vector(to_unsigned(108, 8)),
	122 => std_logic_vector(to_unsigned(106, 8)),
	123 => std_logic_vector(to_unsigned(109, 8)),
	124 => std_logic_vector(to_unsigned(106, 8)),
	125 => std_logic_vector(to_unsigned(109, 8)),
	126 => std_logic_vector(to_unsigned(109, 8)),
	127 => std_logic_vector(to_unsigned(104, 8)),
	128 => std_logic_vector(to_unsigned(103, 8)),
	129 => std_logic_vector(to_unsigned(102, 8)),
	130 => std_logic_vector(to_unsigned(111, 8)),
	131 => std_logic_vector(to_unsigned(103, 8)),
	132 => std_logic_vector(to_unsigned(109, 8)),
	133 => std_logic_vector(to_unsigned(107, 8)),
	134 => std_logic_vector(to_unsigned(107, 8)),
	135 => std_logic_vector(to_unsigned(108, 8)),
	136 => std_logic_vector(to_unsigned(107, 8)),
	137 => std_logic_vector(to_unsigned(110, 8)),
	138 => std_logic_vector(to_unsigned(108, 8)),
	139 => std_logic_vector(to_unsigned(102, 8)),
	140 => std_logic_vector(to_unsigned(103, 8)),
	141 => std_logic_vector(to_unsigned(100, 8)),
	142 => std_logic_vector(to_unsigned(102, 8)),
	143 => std_logic_vector(to_unsigned(110, 8)),
	144 => std_logic_vector(to_unsigned(106, 8)),
	145 => std_logic_vector(to_unsigned(111, 8)),
	146 => std_logic_vector(to_unsigned(107, 8)),
	147 => std_logic_vector(to_unsigned(112, 8)),
	148 => std_logic_vector(to_unsigned(111, 8)),
	149 => std_logic_vector(to_unsigned(105, 8)),
	150 => std_logic_vector(to_unsigned(100, 8)),
	151 => std_logic_vector(to_unsigned(109, 8)),
	152 => std_logic_vector(to_unsigned(109, 8)),
	153 => std_logic_vector(to_unsigned(107, 8)),
	154 => std_logic_vector(to_unsigned(104, 8)),
	155 => std_logic_vector(to_unsigned(106, 8)),
	156 => std_logic_vector(to_unsigned(102, 8)),
	157 => std_logic_vector(to_unsigned(106, 8)),
	158 => std_logic_vector(to_unsigned(104, 8)),
	159 => std_logic_vector(to_unsigned(108, 8)),
	160 => std_logic_vector(to_unsigned(105, 8)),
	161 => std_logic_vector(to_unsigned(104, 8)),
	162 => std_logic_vector(to_unsigned(103, 8)),
	163 => std_logic_vector(to_unsigned(101, 8)),
	164 => std_logic_vector(to_unsigned(106, 8)),
	165 => std_logic_vector(to_unsigned(106, 8)),
	166 => std_logic_vector(to_unsigned(105, 8)),
	167 => std_logic_vector(to_unsigned(103, 8)),
	168 => std_logic_vector(to_unsigned(106, 8)),
	169 => std_logic_vector(to_unsigned(110, 8)),
	170 => std_logic_vector(to_unsigned(111, 8)),
	171 => std_logic_vector(to_unsigned(106, 8)),
	172 => std_logic_vector(to_unsigned(101, 8)),
	173 => std_logic_vector(to_unsigned(112, 8)),
	174 => std_logic_vector(to_unsigned(99, 8)),
	175 => std_logic_vector(to_unsigned(99, 8)),
	176 => std_logic_vector(to_unsigned(106, 8)),
	177 => std_logic_vector(to_unsigned(102, 8)),
	178 => std_logic_vector(to_unsigned(105, 8)),
	179 => std_logic_vector(to_unsigned(106, 8)),
	180 => std_logic_vector(to_unsigned(106, 8)),
	181 => std_logic_vector(to_unsigned(111, 8)),
	182 => std_logic_vector(to_unsigned(106, 8)),
	183 => std_logic_vector(to_unsigned(101, 8)),
	184 => std_logic_vector(to_unsigned(110, 8)),
	185 => std_logic_vector(to_unsigned(110, 8)),
	186 => std_logic_vector(to_unsigned(109, 8)),
	187 => std_logic_vector(to_unsigned(108, 8)),
	188 => std_logic_vector(to_unsigned(100, 8)),
	189 => std_logic_vector(to_unsigned(105, 8)),
	190 => std_logic_vector(to_unsigned(108, 8)),
	191 => std_logic_vector(to_unsigned(107, 8)),
	192 => std_logic_vector(to_unsigned(106, 8)),
	193 => std_logic_vector(to_unsigned(101, 8)),
	194 => std_logic_vector(to_unsigned(104, 8)),
	195 => std_logic_vector(to_unsigned(101, 8)),
	196 => std_logic_vector(to_unsigned(99, 8)),
	197 => std_logic_vector(to_unsigned(109, 8)),
	198 => std_logic_vector(to_unsigned(112, 8)),
	199 => std_logic_vector(to_unsigned(105, 8)),
	200 => std_logic_vector(to_unsigned(105, 8)),
	201 => std_logic_vector(to_unsigned(99, 8)),
	202 => std_logic_vector(to_unsigned(105, 8)),
	203 => std_logic_vector(to_unsigned(99, 8)),
	204 => std_logic_vector(to_unsigned(100, 8)),
	205 => std_logic_vector(to_unsigned(100, 8)),
	206 => std_logic_vector(to_unsigned(100, 8)),
	207 => std_logic_vector(to_unsigned(103, 8)),
	208 => std_logic_vector(to_unsigned(108, 8)),
	209 => std_logic_vector(to_unsigned(111, 8)),
	210 => std_logic_vector(to_unsigned(111, 8)),
	211 => std_logic_vector(to_unsigned(102, 8)),
	212 => std_logic_vector(to_unsigned(104, 8)),
	213 => std_logic_vector(to_unsigned(112, 8)),
	214 => std_logic_vector(to_unsigned(102, 8)),
	215 => std_logic_vector(to_unsigned(106, 8)),
	216 => std_logic_vector(to_unsigned(100, 8)),
	217 => std_logic_vector(to_unsigned(112, 8)),
	218 => std_logic_vector(to_unsigned(100, 8)),
	219 => std_logic_vector(to_unsigned(112, 8)),
	220 => std_logic_vector(to_unsigned(100, 8)),
	221 => std_logic_vector(to_unsigned(99, 8)),
	222 => std_logic_vector(to_unsigned(102, 8)),
	223 => std_logic_vector(to_unsigned(101, 8)),
	224 => std_logic_vector(to_unsigned(100, 8)),
	225 => std_logic_vector(to_unsigned(100, 8)),
	226 => std_logic_vector(to_unsigned(104, 8)),
	227 => std_logic_vector(to_unsigned(106, 8)),
	228 => std_logic_vector(to_unsigned(108, 8)),
	229 => std_logic_vector(to_unsigned(107, 8)),
	230 => std_logic_vector(to_unsigned(101, 8)),
	231 => std_logic_vector(to_unsigned(105, 8)),
	232 => std_logic_vector(to_unsigned(105, 8)),
	233 => std_logic_vector(to_unsigned(101, 8)),
	234 => std_logic_vector(to_unsigned(104, 8)),
	235 => std_logic_vector(to_unsigned(106, 8)),
	236 => std_logic_vector(to_unsigned(105, 8)),
	237 => std_logic_vector(to_unsigned(109, 8)),
	238 => std_logic_vector(to_unsigned(109, 8)),
	239 => std_logic_vector(to_unsigned(112, 8)),
	240 => std_logic_vector(to_unsigned(111, 8)),
	241 => std_logic_vector(to_unsigned(111, 8)),
	242 => std_logic_vector(to_unsigned(111, 8)),
	243 => std_logic_vector(to_unsigned(109, 8)),
	244 => std_logic_vector(to_unsigned(99, 8)),
	245 => std_logic_vector(to_unsigned(102, 8)),
	246 => std_logic_vector(to_unsigned(112, 8)),
	247 => std_logic_vector(to_unsigned(104, 8)),
	248 => std_logic_vector(to_unsigned(107, 8)),
	249 => std_logic_vector(to_unsigned(109, 8)),
	250 => std_logic_vector(to_unsigned(105, 8)),
	251 => std_logic_vector(to_unsigned(103, 8)),
	252 => std_logic_vector(to_unsigned(112, 8)),
	253 => std_logic_vector(to_unsigned(109, 8)),
	254 => std_logic_vector(to_unsigned(109, 8)),
	255 => std_logic_vector(to_unsigned(100, 8)),
	256 => std_logic_vector(to_unsigned(103, 8)),
	257 => std_logic_vector(to_unsigned(106, 8)),
	258 => std_logic_vector(to_unsigned(101, 8)),
	259 => std_logic_vector(to_unsigned(103, 8)),
	260 => std_logic_vector(to_unsigned(106, 8)),
	261 => std_logic_vector(to_unsigned(103, 8)),
	262 => std_logic_vector(to_unsigned(99, 8)),
	263 => std_logic_vector(to_unsigned(104, 8)),
	264 => std_logic_vector(to_unsigned(99, 8)),
	265 => std_logic_vector(to_unsigned(109, 8)),
	266 => std_logic_vector(to_unsigned(107, 8)),
	267 => std_logic_vector(to_unsigned(107, 8)),
	268 => std_logic_vector(to_unsigned(109, 8)),
	269 => std_logic_vector(to_unsigned(106, 8)),
	270 => std_logic_vector(to_unsigned(108, 8)),
	271 => std_logic_vector(to_unsigned(99, 8)),
	272 => std_logic_vector(to_unsigned(103, 8)),
	273 => std_logic_vector(to_unsigned(106, 8)),
	274 => std_logic_vector(to_unsigned(105, 8)),
	275 => std_logic_vector(to_unsigned(107, 8)),
	276 => std_logic_vector(to_unsigned(101, 8)),
	277 => std_logic_vector(to_unsigned(103, 8)),
	278 => std_logic_vector(to_unsigned(109, 8)),
	279 => std_logic_vector(to_unsigned(107, 8)),
	280 => std_logic_vector(to_unsigned(112, 8)),
	281 => std_logic_vector(to_unsigned(109, 8)),
	282 => std_logic_vector(to_unsigned(109, 8)),
	283 => std_logic_vector(to_unsigned(111, 8)),
	284 => std_logic_vector(to_unsigned(106, 8)),
	285 => std_logic_vector(to_unsigned(104, 8)),
	286 => std_logic_vector(to_unsigned(103, 8)),
	287 => std_logic_vector(to_unsigned(103, 8)),
	288 => std_logic_vector(to_unsigned(100, 8)),
	289 => std_logic_vector(to_unsigned(111, 8)),
	290 => std_logic_vector(to_unsigned(107, 8)),
	291 => std_logic_vector(to_unsigned(111, 8)),
	292 => std_logic_vector(to_unsigned(105, 8)),
	293 => std_logic_vector(to_unsigned(109, 8)),
	294 => std_logic_vector(to_unsigned(109, 8)),
	295 => std_logic_vector(to_unsigned(101, 8)),
	296 => std_logic_vector(to_unsigned(108, 8)),
	297 => std_logic_vector(to_unsigned(100, 8)),
	298 => std_logic_vector(to_unsigned(112, 8)),
	299 => std_logic_vector(to_unsigned(108, 8)),
	300 => std_logic_vector(to_unsigned(107, 8)),
	301 => std_logic_vector(to_unsigned(111, 8)),
	302 => std_logic_vector(to_unsigned(111, 8)),
	303 => std_logic_vector(to_unsigned(104, 8)),
	304 => std_logic_vector(to_unsigned(102, 8)),
	305 => std_logic_vector(to_unsigned(103, 8)),
	306 => std_logic_vector(to_unsigned(103, 8)),
	307 => std_logic_vector(to_unsigned(110, 8)),
	308 => std_logic_vector(to_unsigned(100, 8)),
	309 => std_logic_vector(to_unsigned(99, 8)),
	310 => std_logic_vector(to_unsigned(101, 8)),
	311 => std_logic_vector(to_unsigned(100, 8)),
	312 => std_logic_vector(to_unsigned(112, 8)),
	313 => std_logic_vector(to_unsigned(108, 8)),
	314 => std_logic_vector(to_unsigned(111, 8)),
	315 => std_logic_vector(to_unsigned(105, 8)),
	316 => std_logic_vector(to_unsigned(103, 8)),
	317 => std_logic_vector(to_unsigned(107, 8)),
	318 => std_logic_vector(to_unsigned(101, 8)),
	319 => std_logic_vector(to_unsigned(107, 8)),
	320 => std_logic_vector(to_unsigned(105, 8)),
	321 => std_logic_vector(to_unsigned(102, 8)),
	322 => std_logic_vector(to_unsigned(106, 8)),
	323 => std_logic_vector(to_unsigned(99, 8)),
	324 => std_logic_vector(to_unsigned(103, 8)),
	325 => std_logic_vector(to_unsigned(107, 8)),
	326 => std_logic_vector(to_unsigned(109, 8)),
	327 => std_logic_vector(to_unsigned(104, 8)),
	328 => std_logic_vector(to_unsigned(106, 8)),
	329 => std_logic_vector(to_unsigned(106, 8)),
	330 => std_logic_vector(to_unsigned(99, 8)),
	331 => std_logic_vector(to_unsigned(102, 8)),
	332 => std_logic_vector(to_unsigned(100, 8)),
	333 => std_logic_vector(to_unsigned(103, 8)),
	334 => std_logic_vector(to_unsigned(112, 8)),
	335 => std_logic_vector(to_unsigned(110, 8)),
	336 => std_logic_vector(to_unsigned(106, 8)),
	337 => std_logic_vector(to_unsigned(109, 8)),
	338 => std_logic_vector(to_unsigned(100, 8)),
	339 => std_logic_vector(to_unsigned(100, 8)),
	340 => std_logic_vector(to_unsigned(103, 8)),
	341 => std_logic_vector(to_unsigned(102, 8)),
	342 => std_logic_vector(to_unsigned(106, 8)),
	343 => std_logic_vector(to_unsigned(112, 8)),
	344 => std_logic_vector(to_unsigned(104, 8)),
	345 => std_logic_vector(to_unsigned(112, 8)),
	346 => std_logic_vector(to_unsigned(112, 8)),
	347 => std_logic_vector(to_unsigned(110, 8)),
	348 => std_logic_vector(to_unsigned(111, 8)),
	349 => std_logic_vector(to_unsigned(112, 8)),
	350 => std_logic_vector(to_unsigned(112, 8)),
	351 => std_logic_vector(to_unsigned(112, 8)),
	352 => std_logic_vector(to_unsigned(101, 8)),
	353 => std_logic_vector(to_unsigned(105, 8)),
	354 => std_logic_vector(to_unsigned(100, 8)),
	355 => std_logic_vector(to_unsigned(106, 8)),
	356 => std_logic_vector(to_unsigned(106, 8)),
	357 => std_logic_vector(to_unsigned(105, 8)),
	358 => std_logic_vector(to_unsigned(111, 8)),
	359 => std_logic_vector(to_unsigned(110, 8)),
	360 => std_logic_vector(to_unsigned(111, 8)),
	361 => std_logic_vector(to_unsigned(102, 8)),
	362 => std_logic_vector(to_unsigned(106, 8)),
	363 => std_logic_vector(to_unsigned(110, 8)),
	364 => std_logic_vector(to_unsigned(106, 8)),
	365 => std_logic_vector(to_unsigned(103, 8)),
	366 => std_logic_vector(to_unsigned(108, 8)),
	367 => std_logic_vector(to_unsigned(109, 8)),
	368 => std_logic_vector(to_unsigned(106, 8)),
	369 => std_logic_vector(to_unsigned(105, 8)),
	370 => std_logic_vector(to_unsigned(112, 8)),
	371 => std_logic_vector(to_unsigned(104, 8)),
	372 => std_logic_vector(to_unsigned(109, 8)),
	373 => std_logic_vector(to_unsigned(110, 8)),
	374 => std_logic_vector(to_unsigned(99, 8)),
	375 => std_logic_vector(to_unsigned(104, 8)),
	376 => std_logic_vector(to_unsigned(111, 8)),
	377 => std_logic_vector(to_unsigned(110, 8)),
	378 => std_logic_vector(to_unsigned(110, 8)),
	379 => std_logic_vector(to_unsigned(102, 8)),
	380 => std_logic_vector(to_unsigned(105, 8)),
	381 => std_logic_vector(to_unsigned(106, 8)),
	382 => std_logic_vector(to_unsigned(106, 8)),
	others =>(others =>'0'));

component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_rst         : in  std_logic;
      i_start       : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector (7 downto 0)
      );
end component project_reti_logiche;


begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_rst      	=> tb_rst,
          i_start       => tb_start,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
          o_we 		=> mem_we,
          o_data    	=> mem_i_data
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;


MEM : process(tb_clk, tb_start)
begin
    if tb_clk'event and tb_clk = '1' then
        if enable_wire = '1' then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
            end if;
        end if;
    end if;
		if (rising_edge(tb_start)) then
			if (RAM(763) = std_logic_vector(to_unsigned(224, 8))) then
				RAM <= (0 => std_logic_vector(to_unsigned(2, 8)),
		    	1 => std_logic_vector(to_unsigned(12, 8)),
		    	2 => std_logic_vector(to_unsigned(54, 8)),
		    	3 => std_logic_vector(to_unsigned(32, 8)),
		    	4 => std_logic_vector(to_unsigned(50, 8)),
		    	5 => std_logic_vector(to_unsigned(25, 8)),
		    	6 => std_logic_vector(to_unsigned(39, 8)),
		    	7 => std_logic_vector(to_unsigned(70, 8)),
		    	8 => std_logic_vector(to_unsigned(56, 8)),
		    	9 => std_logic_vector(to_unsigned(72, 8)),
		    	10 => std_logic_vector(to_unsigned(73, 8)),
		    	11 => std_logic_vector(to_unsigned(41, 8)),
		    	12 => std_logic_vector(to_unsigned(75, 8)),
		    	13 => std_logic_vector(to_unsigned(72, 8)),
		    	14 => std_logic_vector(to_unsigned(32, 8)),
		    	15 => std_logic_vector(to_unsigned(67, 8)),
		    	16 => std_logic_vector(to_unsigned(58, 8)),
		    	17 => std_logic_vector(to_unsigned(47, 8)),
		    	18 => std_logic_vector(to_unsigned(39, 8)),
		    	19 => std_logic_vector(to_unsigned(28, 8)),
		    	20 => std_logic_vector(to_unsigned(65, 8)),
		    	21 => std_logic_vector(to_unsigned(75, 8)),
		    	22 => std_logic_vector(to_unsigned(71, 8)),
		    	23 => std_logic_vector(to_unsigned(62, 8)),
		    	24 => std_logic_vector(to_unsigned(38, 8)),
		    	25 => std_logic_vector(to_unsigned(63, 8)),
		    	others =>(others =>'0'));
			end if;
		end if;
end process;


test : process is
begin
    wait for 100 ns;
    wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_rst <= '0';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;

		assert RAM(383) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(383)))) severity failure;
		assert RAM(384) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(384)))) severity failure;
		assert RAM(385) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(385)))) severity failure;
		assert RAM(386) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(386)))) severity failure;
		assert RAM(387) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(387)))) severity failure;
		assert RAM(388) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(388)))) severity failure;
		assert RAM(389) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(389)))) severity failure;
		assert RAM(390) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(390)))) severity failure;
		assert RAM(391) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(391)))) severity failure;
		assert RAM(392) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(392)))) severity failure;
		assert RAM(393) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(393)))) severity failure;
		assert RAM(394) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(394)))) severity failure;
		assert RAM(395) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(395)))) severity failure;
		assert RAM(396) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(396)))) severity failure;
		assert RAM(397) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(397)))) severity failure;
		assert RAM(398) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(398)))) severity failure;
		assert RAM(399) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(399)))) severity failure;
		assert RAM(400) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(400)))) severity failure;
		assert RAM(401) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(401)))) severity failure;
		assert RAM(402) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(402)))) severity failure;
		assert RAM(403) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(403)))) severity failure;
		assert RAM(404) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(404)))) severity failure;
		assert RAM(405) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(405)))) severity failure;
		assert RAM(406) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(406)))) severity failure;
		assert RAM(407) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(407)))) severity failure;
		assert RAM(408) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(408)))) severity failure;
		assert RAM(409) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(409)))) severity failure;
		assert RAM(410) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(410)))) severity failure;
		assert RAM(411) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(411)))) severity failure;
		assert RAM(412) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(412)))) severity failure;
		assert RAM(413) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(413)))) severity failure;
		assert RAM(414) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(414)))) severity failure;
		assert RAM(415) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(415)))) severity failure;
		assert RAM(416) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(416)))) severity failure;
		assert RAM(417) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(417)))) severity failure;
		assert RAM(418) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(418)))) severity failure;
		assert RAM(419) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(419)))) severity failure;
		assert RAM(420) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(420)))) severity failure;
		assert RAM(421) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(421)))) severity failure;
		assert RAM(422) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(422)))) severity failure;
		assert RAM(423) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(423)))) severity failure;
		assert RAM(424) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(424)))) severity failure;
		assert RAM(425) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(425)))) severity failure;
		assert RAM(426) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(426)))) severity failure;
		assert RAM(427) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(427)))) severity failure;
		assert RAM(428) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(428)))) severity failure;
		assert RAM(429) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(429)))) severity failure;
		assert RAM(430) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(430)))) severity failure;
		assert RAM(431) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(431)))) severity failure;
		assert RAM(432) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(432)))) severity failure;
		assert RAM(433) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(433)))) severity failure;
		assert RAM(434) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(434)))) severity failure;
		assert RAM(435) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(435)))) severity failure;
		assert RAM(436) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(436)))) severity failure;
		assert RAM(437) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(437)))) severity failure;
		assert RAM(438) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(438)))) severity failure;
		assert RAM(439) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(439)))) severity failure;
		assert RAM(440) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(440)))) severity failure;
		assert RAM(441) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(441)))) severity failure;
		assert RAM(442) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(442)))) severity failure;
		assert RAM(443) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(443)))) severity failure;
		assert RAM(444) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(444)))) severity failure;
		assert RAM(445) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(445)))) severity failure;
		assert RAM(446) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(446)))) severity failure;
		assert RAM(447) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(447)))) severity failure;
		assert RAM(448) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(448)))) severity failure;
		assert RAM(449) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(449)))) severity failure;
		assert RAM(450) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(450)))) severity failure;
		assert RAM(451) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(451)))) severity failure;
		assert RAM(452) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(452)))) severity failure;
		assert RAM(453) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(453)))) severity failure;
		assert RAM(454) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(454)))) severity failure;
		assert RAM(455) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(455)))) severity failure;
		assert RAM(456) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(456)))) severity failure;
		assert RAM(457) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(457)))) severity failure;
		assert RAM(458) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(458)))) severity failure;
		assert RAM(459) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(459)))) severity failure;
		assert RAM(460) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(460)))) severity failure;
		assert RAM(461) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(461)))) severity failure;
		assert RAM(462) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(462)))) severity failure;
		assert RAM(463) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(463)))) severity failure;
		assert RAM(464) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(464)))) severity failure;
		assert RAM(465) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(465)))) severity failure;
		assert RAM(466) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(466)))) severity failure;
		assert RAM(467) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(467)))) severity failure;
		assert RAM(468) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(468)))) severity failure;
		assert RAM(469) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(469)))) severity failure;
		assert RAM(470) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(470)))) severity failure;
		assert RAM(471) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(471)))) severity failure;
		assert RAM(472) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(472)))) severity failure;
		assert RAM(473) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(473)))) severity failure;
		assert RAM(474) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(474)))) severity failure;
		assert RAM(475) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(475)))) severity failure;
		assert RAM(476) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(476)))) severity failure;
		assert RAM(477) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(477)))) severity failure;
		assert RAM(478) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(478)))) severity failure;
		assert RAM(479) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(479)))) severity failure;
		assert RAM(480) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(480)))) severity failure;
		assert RAM(481) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(481)))) severity failure;
		assert RAM(482) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(482)))) severity failure;
		assert RAM(483) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(483)))) severity failure;
		assert RAM(484) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(484)))) severity failure;
		assert RAM(485) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(485)))) severity failure;
		assert RAM(486) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(486)))) severity failure;
		assert RAM(487) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(487)))) severity failure;
		assert RAM(488) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(488)))) severity failure;
		assert RAM(489) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(489)))) severity failure;
		assert RAM(490) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(490)))) severity failure;
		assert RAM(491) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(491)))) severity failure;
		assert RAM(492) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(492)))) severity failure;
		assert RAM(493) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(493)))) severity failure;
		assert RAM(494) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(494)))) severity failure;
		assert RAM(495) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(495)))) severity failure;
		assert RAM(496) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(496)))) severity failure;
		assert RAM(497) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(497)))) severity failure;
		assert RAM(498) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(498)))) severity failure;
		assert RAM(499) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(499)))) severity failure;
		assert RAM(500) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(500)))) severity failure;
		assert RAM(501) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(501)))) severity failure;
		assert RAM(502) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(502)))) severity failure;
		assert RAM(503) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(503)))) severity failure;
		assert RAM(504) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(504)))) severity failure;
		assert RAM(505) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(505)))) severity failure;
		assert RAM(506) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(506)))) severity failure;
		assert RAM(507) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(507)))) severity failure;
		assert RAM(508) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(508)))) severity failure;
		assert RAM(509) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(509)))) severity failure;
		assert RAM(510) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(510)))) severity failure;
		assert RAM(511) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(511)))) severity failure;
		assert RAM(512) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(512)))) severity failure;
		assert RAM(513) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(513)))) severity failure;
		assert RAM(514) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(514)))) severity failure;
		assert RAM(515) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(515)))) severity failure;
		assert RAM(516) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(516)))) severity failure;
		assert RAM(517) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(517)))) severity failure;
		assert RAM(518) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(518)))) severity failure;
		assert RAM(519) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(519)))) severity failure;
		assert RAM(520) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(520)))) severity failure;
		assert RAM(521) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(521)))) severity failure;
		assert RAM(522) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(522)))) severity failure;
		assert RAM(523) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(523)))) severity failure;
		assert RAM(524) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(524)))) severity failure;
		assert RAM(525) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(525)))) severity failure;
		assert RAM(526) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(526)))) severity failure;
		assert RAM(527) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(527)))) severity failure;
		assert RAM(528) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(528)))) severity failure;
		assert RAM(529) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(529)))) severity failure;
		assert RAM(530) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(530)))) severity failure;
		assert RAM(531) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(531)))) severity failure;
		assert RAM(532) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(532)))) severity failure;
		assert RAM(533) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(533)))) severity failure;
		assert RAM(534) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(534)))) severity failure;
		assert RAM(535) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(535)))) severity failure;
		assert RAM(536) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(536)))) severity failure;
		assert RAM(537) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(537)))) severity failure;
		assert RAM(538) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(538)))) severity failure;
		assert RAM(539) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(539)))) severity failure;
		assert RAM(540) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(540)))) severity failure;
		assert RAM(541) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(541)))) severity failure;
		assert RAM(542) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(542)))) severity failure;
		assert RAM(543) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(543)))) severity failure;
		assert RAM(544) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(544)))) severity failure;
		assert RAM(545) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(545)))) severity failure;
		assert RAM(546) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(546)))) severity failure;
		assert RAM(547) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(547)))) severity failure;
		assert RAM(548) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(548)))) severity failure;
		assert RAM(549) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(549)))) severity failure;
		assert RAM(550) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(550)))) severity failure;
		assert RAM(551) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(551)))) severity failure;
		assert RAM(552) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(552)))) severity failure;
		assert RAM(553) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(553)))) severity failure;
		assert RAM(554) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(554)))) severity failure;
		assert RAM(555) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(555)))) severity failure;
		assert RAM(556) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(556)))) severity failure;
		assert RAM(557) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(557)))) severity failure;
		assert RAM(558) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(558)))) severity failure;
		assert RAM(559) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(559)))) severity failure;
		assert RAM(560) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(560)))) severity failure;
		assert RAM(561) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(561)))) severity failure;
		assert RAM(562) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(562)))) severity failure;
		assert RAM(563) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(563)))) severity failure;
		assert RAM(564) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(564)))) severity failure;
		assert RAM(565) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(565)))) severity failure;
		assert RAM(566) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(566)))) severity failure;
		assert RAM(567) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(567)))) severity failure;
		assert RAM(568) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(568)))) severity failure;
		assert RAM(569) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(569)))) severity failure;
		assert RAM(570) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(570)))) severity failure;
		assert RAM(571) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(571)))) severity failure;
		assert RAM(572) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(572)))) severity failure;
		assert RAM(573) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(573)))) severity failure;
		assert RAM(574) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(574)))) severity failure;
		assert RAM(575) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(575)))) severity failure;
		assert RAM(576) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(576)))) severity failure;
		assert RAM(577) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(577)))) severity failure;
		assert RAM(578) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(578)))) severity failure;
		assert RAM(579) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(579)))) severity failure;
		assert RAM(580) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(580)))) severity failure;
		assert RAM(581) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(581)))) severity failure;
		assert RAM(582) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(582)))) severity failure;
		assert RAM(583) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(583)))) severity failure;
		assert RAM(584) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(584)))) severity failure;
		assert RAM(585) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(585)))) severity failure;
		assert RAM(586) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(586)))) severity failure;
		assert RAM(587) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(587)))) severity failure;
		assert RAM(588) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(588)))) severity failure;
		assert RAM(589) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(589)))) severity failure;
		assert RAM(590) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(590)))) severity failure;
		assert RAM(591) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(591)))) severity failure;
		assert RAM(592) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(592)))) severity failure;
		assert RAM(593) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(593)))) severity failure;
		assert RAM(594) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(594)))) severity failure;
		assert RAM(595) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(595)))) severity failure;
		assert RAM(596) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(596)))) severity failure;
		assert RAM(597) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(597)))) severity failure;
		assert RAM(598) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(598)))) severity failure;
		assert RAM(599) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(599)))) severity failure;
		assert RAM(600) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(600)))) severity failure;
		assert RAM(601) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(601)))) severity failure;
		assert RAM(602) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(602)))) severity failure;
		assert RAM(603) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(603)))) severity failure;
		assert RAM(604) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(604)))) severity failure;
		assert RAM(605) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(605)))) severity failure;
		assert RAM(606) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(606)))) severity failure;
		assert RAM(607) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(607)))) severity failure;
		assert RAM(608) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(608)))) severity failure;
		assert RAM(609) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(609)))) severity failure;
		assert RAM(610) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(610)))) severity failure;
		assert RAM(611) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(611)))) severity failure;
		assert RAM(612) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(612)))) severity failure;
		assert RAM(613) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(613)))) severity failure;
		assert RAM(614) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(614)))) severity failure;
		assert RAM(615) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(615)))) severity failure;
		assert RAM(616) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(616)))) severity failure;
		assert RAM(617) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(617)))) severity failure;
		assert RAM(618) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(618)))) severity failure;
		assert RAM(619) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(619)))) severity failure;
		assert RAM(620) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(620)))) severity failure;
		assert RAM(621) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(621)))) severity failure;
		assert RAM(622) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(622)))) severity failure;
		assert RAM(623) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(623)))) severity failure;
		assert RAM(624) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(624)))) severity failure;
		assert RAM(625) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(625)))) severity failure;
		assert RAM(626) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(626)))) severity failure;
		assert RAM(627) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(627)))) severity failure;
		assert RAM(628) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(628)))) severity failure;
		assert RAM(629) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(629)))) severity failure;
		assert RAM(630) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(630)))) severity failure;
		assert RAM(631) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(631)))) severity failure;
		assert RAM(632) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(632)))) severity failure;
		assert RAM(633) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(633)))) severity failure;
		assert RAM(634) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(634)))) severity failure;
		assert RAM(635) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(635)))) severity failure;
		assert RAM(636) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(636)))) severity failure;
		assert RAM(637) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(637)))) severity failure;
		assert RAM(638) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(638)))) severity failure;
		assert RAM(639) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(639)))) severity failure;
		assert RAM(640) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(640)))) severity failure;
		assert RAM(641) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(641)))) severity failure;
		assert RAM(642) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(642)))) severity failure;
		assert RAM(643) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(643)))) severity failure;
		assert RAM(644) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(644)))) severity failure;
		assert RAM(645) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(645)))) severity failure;
		assert RAM(646) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(646)))) severity failure;
		assert RAM(647) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(647)))) severity failure;
		assert RAM(648) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(648)))) severity failure;
		assert RAM(649) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(649)))) severity failure;
		assert RAM(650) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(650)))) severity failure;
		assert RAM(651) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(651)))) severity failure;
		assert RAM(652) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(652)))) severity failure;
		assert RAM(653) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(653)))) severity failure;
		assert RAM(654) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(654)))) severity failure;
		assert RAM(655) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(655)))) severity failure;
		assert RAM(656) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(656)))) severity failure;
		assert RAM(657) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(657)))) severity failure;
		assert RAM(658) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(658)))) severity failure;
		assert RAM(659) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(659)))) severity failure;
		assert RAM(660) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(660)))) severity failure;
		assert RAM(661) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(661)))) severity failure;
		assert RAM(662) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(662)))) severity failure;
		assert RAM(663) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(663)))) severity failure;
		assert RAM(664) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(664)))) severity failure;
		assert RAM(665) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(665)))) severity failure;
		assert RAM(666) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(666)))) severity failure;
		assert RAM(667) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(667)))) severity failure;
		assert RAM(668) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(668)))) severity failure;
		assert RAM(669) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(669)))) severity failure;
		assert RAM(670) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(670)))) severity failure;
		assert RAM(671) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(671)))) severity failure;
		assert RAM(672) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(672)))) severity failure;
		assert RAM(673) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(673)))) severity failure;
		assert RAM(674) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(674)))) severity failure;
		assert RAM(675) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(675)))) severity failure;
		assert RAM(676) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(676)))) severity failure;
		assert RAM(677) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(677)))) severity failure;
		assert RAM(678) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(678)))) severity failure;
		assert RAM(679) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(679)))) severity failure;
		assert RAM(680) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(680)))) severity failure;
		assert RAM(681) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(681)))) severity failure;
		assert RAM(682) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(682)))) severity failure;
		assert RAM(683) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(683)))) severity failure;
		assert RAM(684) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(684)))) severity failure;
		assert RAM(685) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(685)))) severity failure;
		assert RAM(686) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(686)))) severity failure;
		assert RAM(687) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(687)))) severity failure;
		assert RAM(688) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(688)))) severity failure;
		assert RAM(689) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(689)))) severity failure;
		assert RAM(690) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(690)))) severity failure;
		assert RAM(691) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(691)))) severity failure;
		assert RAM(692) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(692)))) severity failure;
		assert RAM(693) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(693)))) severity failure;
		assert RAM(694) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(694)))) severity failure;
		assert RAM(695) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(695)))) severity failure;
		assert RAM(696) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(696)))) severity failure;
		assert RAM(697) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(697)))) severity failure;
		assert RAM(698) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(698)))) severity failure;
		assert RAM(699) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(699)))) severity failure;
		assert RAM(700) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(700)))) severity failure;
		assert RAM(701) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(701)))) severity failure;
		assert RAM(702) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(702)))) severity failure;
		assert RAM(703) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(703)))) severity failure;
		assert RAM(704) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(704)))) severity failure;
		assert RAM(705) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(705)))) severity failure;
		assert RAM(706) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(706)))) severity failure;
		assert RAM(707) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(707)))) severity failure;
		assert RAM(708) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(708)))) severity failure;
		assert RAM(709) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(709)))) severity failure;
		assert RAM(710) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(710)))) severity failure;
		assert RAM(711) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(711)))) severity failure;
		assert RAM(712) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(712)))) severity failure;
		assert RAM(713) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(713)))) severity failure;
		assert RAM(714) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(714)))) severity failure;
		assert RAM(715) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(715)))) severity failure;
		assert RAM(716) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(716)))) severity failure;
		assert RAM(717) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(717)))) severity failure;
		assert RAM(718) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(718)))) severity failure;
		assert RAM(719) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(719)))) severity failure;
		assert RAM(720) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(720)))) severity failure;
		assert RAM(721) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(721)))) severity failure;
		assert RAM(722) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(722)))) severity failure;
		assert RAM(723) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(723)))) severity failure;
		assert RAM(724) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(724)))) severity failure;
		assert RAM(725) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(725)))) severity failure;
		assert RAM(726) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(726)))) severity failure;
		assert RAM(727) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(727)))) severity failure;
		assert RAM(728) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(728)))) severity failure;
		assert RAM(729) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(729)))) severity failure;
		assert RAM(730) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(730)))) severity failure;
		assert RAM(731) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(731)))) severity failure;
		assert RAM(732) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(732)))) severity failure;
		assert RAM(733) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected 64 found " & integer'image(to_integer(unsigned(RAM(733)))) severity failure;
		assert RAM(734) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(734)))) severity failure;
		assert RAM(735) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected 32 found " & integer'image(to_integer(unsigned(RAM(735)))) severity failure;
		assert RAM(736) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(736)))) severity failure;
		assert RAM(737) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(737)))) severity failure;
		assert RAM(738) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(738)))) severity failure;
		assert RAM(739) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(739)))) severity failure;
		assert RAM(740) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(740)))) severity failure;
		assert RAM(741) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(741)))) severity failure;
		assert RAM(742) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(742)))) severity failure;
		assert RAM(743) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(743)))) severity failure;
		assert RAM(744) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(744)))) severity failure;
		assert RAM(745) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(745)))) severity failure;
		assert RAM(746) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(746)))) severity failure;
		assert RAM(747) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(747)))) severity failure;
		assert RAM(748) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(748)))) severity failure;
		assert RAM(749) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(749)))) severity failure;
		assert RAM(750) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(750)))) severity failure;
		assert RAM(751) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(751)))) severity failure;
		assert RAM(752) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(752)))) severity failure;
		assert RAM(753) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(753)))) severity failure;
		assert RAM(754) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(754)))) severity failure;
		assert RAM(755) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(755)))) severity failure;
		assert RAM(756) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected 160 found " & integer'image(to_integer(unsigned(RAM(756)))) severity failure;
		assert RAM(757) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(757)))) severity failure;
		assert RAM(758) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(758)))) severity failure;
		assert RAM(759) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(759)))) severity failure;
		assert RAM(760) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected 96 found " & integer'image(to_integer(unsigned(RAM(760)))) severity failure;
		assert RAM(761) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected 192 found " & integer'image(to_integer(unsigned(RAM(761)))) severity failure;
		assert RAM(762) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(762)))) severity failure;
		assert RAM(763) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected 224 found " & integer'image(to_integer(unsigned(RAM(763)))) severity failure;

		wait for 100 ns;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;

		assert RAM(26) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected 232 found " & integer'image(to_integer(unsigned(RAM(26)))) severity failure;
    assert RAM(27) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected 56 found " & integer'image(to_integer(unsigned(RAM(27)))) severity failure;
    assert RAM(28) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected 200 found " & integer'image(to_integer(unsigned(RAM(28)))) severity failure;
    assert RAM(29) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected 0 found " & integer'image(to_integer(unsigned(RAM(29)))) severity failure;
    assert RAM(30) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(30)))) severity failure;
    assert RAM(31) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(31)))) severity failure;
    assert RAM(32) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected 248 found " & integer'image(to_integer(unsigned(RAM(32)))) severity failure;
    assert RAM(33) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(33)))) severity failure;
    assert RAM(34) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(34)))) severity failure;
    assert RAM(35) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected 128 found " & integer'image(to_integer(unsigned(RAM(35)))) severity failure;
    assert RAM(36) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(36)))) severity failure;
    assert RAM(37) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(37)))) severity failure;
    assert RAM(38) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected 56 found " & integer'image(to_integer(unsigned(RAM(38)))) severity failure;
    assert RAM(39) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(39)))) severity failure;
    assert RAM(40) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(40)))) severity failure;
    assert RAM(41) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected 176 found " & integer'image(to_integer(unsigned(RAM(41)))) severity failure;
    assert RAM(42) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected 112 found " & integer'image(to_integer(unsigned(RAM(42)))) severity failure;
    assert RAM(43) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected 24 found " & integer'image(to_integer(unsigned(RAM(43)))) severity failure;
    assert RAM(44) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(44)))) severity failure;
    assert RAM(45) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(45)))) severity failure;
    assert RAM(46) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(46)))) severity failure;
    assert RAM(47) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(47)))) severity failure;
    assert RAM(48) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected 104 found " & integer'image(to_integer(unsigned(RAM(48)))) severity failure;
    assert RAM(49) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected 255 found " & integer'image(to_integer(unsigned(RAM(49)))) severity failure;

    assert false report "Simulation Ended! TEST PASSATO" severity failure;
end process test;

end consimgtb;
